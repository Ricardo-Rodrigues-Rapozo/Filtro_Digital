module procTest_00 (

input  clk, rst,
input  signed [31:0] in ,
output signed [31:0] out,
output [0:0] req_in,
output [6:0] out_en);

wire itr = 1'b0;
wire proc_req_in, proc_out_en;
wire [0:0] addr_in;
wire [2:0] addr_out;

`ifdef __ICARUS__
wire mem_wr;
wire [10:0] mem_addr_wr;
wire [8:0] pc_sim_val;
`endif

processor#(.NUBITS(32),
.NBMANT(23),
.NBEXPO(8),
.NBOPER(11),
.NUGAIN(128),
.MDATAS(1824),
.MINSTS(324),
.SDEPTH(5),
.DDEPTH(5),
.NBIOIN(1),
.NBIOOU(3),
.FFTSIZ(7),
.CAL(1),
.SET(1),
.LOD(1),
.LES(1),
.JIZ(1),
.MLT(1),
.ADD(1),
.LDI(1),
.P_LOD(1),
.ILI(1),
.SET_P(1),
.F_MLT(1),
.SF_SU2(1),
.SF_ADD(1),
.F_SU1(1),
.ISI(1),
.F_ADD(1),
.NEG_M(1),
.GRE(1),
.P_NEG_M(1),
.STI(1),
.P_INN(1),
.I2F(1),
.SF_DIV(1),
.EQU(1),
.SF_MLT(1),
.P_I2F_M(1),
.POP(1),
.F2I(1),
.OUT(1),
.DFILE("C:/Users/Ricardo/Desktop/Dissertacao/banco_filtro/procTest_00/Hardware/procTest_00_data.mif"),
.IFILE("C:/Users/Ricardo/Desktop/Dissertacao/banco_filtro/procTest_00/Hardware/procTest_00_inst.mif"))

`ifdef __ICARUS__
p_procTest_00 (clk, rst, in, out, addr_in, addr_out, proc_req_in, proc_out_en, itr, mem_wr, mem_addr_wr,pc_sim_val);
`else
p_procTest_00 (clk, rst, in, out, addr_in, addr_out, proc_req_in, proc_out_en, itr);
`endif

assign req_in = proc_req_in;
addr_dec #(7) dec_out(proc_out_en, addr_out, out_en);

// ----------------------------------------------------------------------------
// Simulacao ------------------------------------------------------------------
// ----------------------------------------------------------------------------

`ifdef __ICARUS__

// I/O ------------------------------------------------------------------------

reg signed [31:0] in_sim_0 = 0;
reg req_in_sim_0 = 0;

reg signed [31:0] out_sig_1 = 0;
reg out_en_sim_1 = 0;
reg signed [31:0] out_sig_2 = 0;
reg out_en_sim_2 = 0;
reg signed [31:0] out_sig_3 = 0;
reg out_en_sim_3 = 0;
reg signed [31:0] out_sig_4 = 0;
reg out_en_sim_4 = 0;
reg signed [31:0] out_sig_5 = 0;
reg out_en_sim_5 = 0;
reg signed [31:0] out_sig_6 = 0;
reg out_en_sim_6 = 0;

always @ (*) begin
   if (req_in == 1) in_sim_0 = in;
   req_in_sim_0 = req_in == 1;
end

always @ (*) begin
   if (out_en == 2) out_sig_1 <= out;
   out_en_sim_1 = out_en == 2;
   if (out_en == 4) out_sig_2 <= out;
   out_en_sim_2 = out_en == 4;
   if (out_en == 8) out_sig_3 <= out;
   out_en_sim_3 = out_en == 8;
   if (out_en == 16) out_sig_4 <= out;
   out_en_sim_4 = out_en == 16;
   if (out_en == 32) out_sig_5 <= out;
   out_en_sim_5 = out_en == 32;
   if (out_en == 64) out_sig_6 <= out;
   out_en_sim_6 = out_en == 64;
end

// variaveis ------------------------------------------------------------------

reg [31:0] me1_f_ifft_v_N_e_ = 0;
reg [31:0] me1_f_ifft_v_mmax_e_ = 0;
reg [31:0] me1_f_ifft_v_istep_e_ = 0;
reg [31:0] me1_f_ifft_v_m_e_ = 0;
reg [31:0] me1_f_ifft_v_ind_e_ = 0;
reg [31:0] me1_f_ifft_v_sind_e_ = 0;
reg [31:0] me1_f_ifft_v_k_e_ = 0;
reg [31:0] me1_f_ifft_v_j_e_ = 0;
reg [31:0] me3_f_ifft_v_temp_i_e_ = 31'dx;
reg [31:0] me3_f_ifft_v_temp_e_ = 31'dx;
reg [31:0] me1_f_main_v_sample_count_e_ = 0;
reg [31:0] me1_f_main_v_output_count_e_ = 0;
reg [31:0] me1_f_main_v_M_e_ = 0;
reg [31:0] me1_f_main_v_fft_limit_e_ = 0;
reg [31:0] me1_f_main_v_k_e_ = 0;
reg [31:0] me1_f_main_v_mm_e_ = 0;

always @ (posedge clk) begin
   if (mem_addr_wr == 384 && mem_wr) me1_f_ifft_v_N_e_ <= out;
   if (mem_addr_wr == 386 && mem_wr) me1_f_ifft_v_mmax_e_ <= out;
   if (mem_addr_wr == 388 && mem_wr) me1_f_ifft_v_istep_e_ <= out;
   if (mem_addr_wr == 390 && mem_wr) me1_f_ifft_v_m_e_ <= out;
   if (mem_addr_wr == 391 && mem_wr) me1_f_ifft_v_ind_e_ <= out;
   if (mem_addr_wr == 392 && mem_wr) me1_f_ifft_v_sind_e_ <= out;
   if (mem_addr_wr == 393 && mem_wr) me1_f_ifft_v_k_e_ <= out;
   if (mem_addr_wr == 394 && mem_wr) me1_f_ifft_v_j_e_ <= out;
   if (mem_addr_wr == 399 && mem_wr) me3_f_ifft_v_temp_i_e_ <= out;
   if (mem_addr_wr == 400 && mem_wr) me3_f_ifft_v_temp_e_ <= out;
   if (mem_addr_wr == 401 && mem_wr) me1_f_main_v_sample_count_e_ <= out;
   if (mem_addr_wr == 402 && mem_wr) me1_f_main_v_output_count_e_ <= out;
   if (mem_addr_wr == 1815 && mem_wr) me1_f_main_v_M_e_ <= out;
   if (mem_addr_wr == 1816 && mem_wr) me1_f_main_v_fft_limit_e_ <= out;
   if (mem_addr_wr == 1817 && mem_wr) me1_f_main_v_k_e_ <= out;
   if (mem_addr_wr == 1819 && mem_wr) me1_f_main_v_mm_e_ <= out;
end

wire [16+32*2-1:0] comp_me3_f_ifft_v_temp_e_ = {8'd23, 8'd8, me3_f_ifft_v_temp_e_, me3_f_ifft_v_temp_i_e_};

// arrays ---------------------------------------------------------------------

reg [32-1:0] arr_me3_f_global_v_E0_e_0000=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0001=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0002=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0003=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0004=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0005=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0006=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0007=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0008=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0009=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0010=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0011=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0012=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0013=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0014=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0015=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0016=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0017=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0018=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0019=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0020=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0021=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0022=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0023=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0024=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0025=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0026=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0027=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0028=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0029=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0030=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0031=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0032=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0033=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0034=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0035=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0036=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0037=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0038=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0039=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0040=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0041=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0042=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0043=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0044=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0045=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0046=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0047=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0048=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0049=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0050=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0051=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0052=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0053=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0054=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0055=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0056=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0057=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0058=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0059=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0060=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0061=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0062=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0063=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0064=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0065=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0066=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0067=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0068=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0069=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0070=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0071=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0072=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0073=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0074=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0075=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0076=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0077=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0078=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0079=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0080=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0081=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0082=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0083=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0084=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0085=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0086=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0087=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0088=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0089=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0090=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0091=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0092=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0093=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0094=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0095=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0096=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0097=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0098=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0099=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0100=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0101=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0102=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0103=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0104=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0105=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0106=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0107=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0108=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0109=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0110=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0111=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0112=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0113=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0114=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0115=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0116=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0117=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0118=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0119=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0120=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0121=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0122=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0123=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0124=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0125=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0126=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_e_0127=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0000=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0001=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0002=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0003=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0004=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0005=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0006=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0007=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0008=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0009=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0010=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0011=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0012=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0013=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0014=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0015=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0016=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0017=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0018=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0019=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0020=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0021=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0022=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0023=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0024=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0025=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0026=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0027=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0028=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0029=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0030=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0031=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0032=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0033=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0034=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0035=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0036=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0037=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0038=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0039=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0040=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0041=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0042=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0043=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0044=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0045=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0046=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0047=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0048=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0049=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0050=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0051=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0052=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0053=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0054=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0055=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0056=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0057=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0058=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0059=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0060=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0061=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0062=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0063=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0064=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0065=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0066=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0067=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0068=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0069=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0070=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0071=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0072=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0073=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0074=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0075=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0076=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0077=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0078=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0079=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0080=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0081=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0082=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0083=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0084=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0085=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0086=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0087=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0088=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0089=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0090=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0091=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0092=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0093=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0094=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0095=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0096=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0097=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0098=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0099=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0100=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0101=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0102=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0103=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0104=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0105=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0106=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0107=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0108=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0109=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0110=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0111=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0112=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0113=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0114=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0115=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0116=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0117=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0118=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0119=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0120=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0121=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0122=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0123=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0124=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0125=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0126=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_E0_i_e_0127=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_wpv_e_0000=32'b01110101010000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_wpv_e_0001=32'b01110100111111111101100010001000;
reg [32-1:0] arr_me3_f_global_v_wpv_e_0002=32'b01110100111111110110001000110111;
reg [32-1:0] arr_me3_f_global_v_wpv_e_0003=32'b01110100111111101001110101010110;
reg [32-1:0] arr_me3_f_global_v_wpv_e_0004=32'b01110100111111011000101001011111;
reg [32-1:0] arr_me3_f_global_v_wpv_e_0005=32'b01110100111111000010100111111100;
reg [32-1:0] arr_me3_f_global_v_wpv_e_0006=32'b01110100111110100111110100000110;
reg [32-1:0] arr_me3_f_global_v_wpv_e_0007=32'b01110100111110001000010010000100;
reg [32-1:0] arr_me3_f_global_v_wpv_e_0008=32'b01110100111101100100000110101111;
reg [32-1:0] arr_me3_f_global_v_wpv_e_0009=32'b01110100111100111011010111101100;
reg [32-1:0] arr_me3_f_global_v_wpv_e_0010=32'b01110100111100001110001011001100;
reg [32-1:0] arr_me3_f_global_v_wpv_e_0011=32'b01110100111011011100101000001101;
reg [32-1:0] arr_me3_f_global_v_wpv_e_0012=32'b01110100111010100110110110011001;
reg [32-1:0] arr_me3_f_global_v_wpv_e_0013=32'b01110100111001101100111110000001;
reg [32-1:0] arr_me3_f_global_v_wpv_e_0014=32'b01110100111000101111001000000010;
reg [32-1:0] arr_me3_f_global_v_wpv_e_0015=32'b01110100110111101101011101111101;
reg [32-1:0] arr_me3_f_global_v_wpv_e_0016=32'b01110100110110101000001001111010;
reg [32-1:0] arr_me3_f_global_v_wpv_e_0017=32'b01110100110101011111010110100101;
reg [32-1:0] arr_me3_f_global_v_wpv_e_0018=32'b01110100110100010011001111001101;
reg [32-1:0] arr_me3_f_global_v_wpv_e_0019=32'b01110100110011000011111111100000;
reg [32-1:0] arr_me3_f_global_v_wpv_e_0020=32'b01110100110001110001110011101101;
reg [32-1:0] arr_me3_f_global_v_wpv_e_0021=32'b01110100110000011100111000011111;
reg [32-1:0] arr_me3_f_global_v_wpv_e_0022=32'b01110100011110001010110101110101;
reg [32-1:0] arr_me3_f_global_v_wpv_e_0023=32'b01110100011011010111010001000000;
reg [32-1:0] arr_me3_f_global_v_wpv_e_0024=32'b01110100011000011111011110001011;
reg [32-1:0] arr_me3_f_global_v_wpv_e_0025=32'b01110100010101100011111001101010;
reg [32-1:0] arr_me3_f_global_v_wpv_e_0026=32'b01110100010010100101000000011001;
reg [32-1:0] arr_me3_f_global_v_wpv_e_0027=32'b01110011111111000110011111100110;
reg [32-1:0] arr_me3_f_global_v_wpv_e_0028=32'b01110011111000111110001011100001;
reg [32-1:0] arr_me3_f_global_v_wpv_e_0029=32'b01110011110010110010000001000010;
reg [32-1:0] arr_me3_f_global_v_wpv_e_0030=32'b01110011011001000101111010011011;
reg [32-1:0] arr_me3_f_global_v_wpv_e_0031=32'b01110010111001000111110110011000;
reg [32-1:0] arr_me3_f_global_v_wpv_e_0032=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_wpv_e_0033=32'b11110010111001000111110110011000;
reg [32-1:0] arr_me3_f_global_v_wpv_e_0034=32'b11110011011001000101111010011011;
reg [32-1:0] arr_me3_f_global_v_wpv_e_0035=32'b11110011110010110010000001000010;
reg [32-1:0] arr_me3_f_global_v_wpv_e_0036=32'b11110011111000111110001011100001;
reg [32-1:0] arr_me3_f_global_v_wpv_e_0037=32'b11110011111111000110011111100110;
reg [32-1:0] arr_me3_f_global_v_wpv_e_0038=32'b11110100010010100101000000011001;
reg [32-1:0] arr_me3_f_global_v_wpv_e_0039=32'b11110100010101100011111001101010;
reg [32-1:0] arr_me3_f_global_v_wpv_e_0040=32'b11110100011000011111011110001011;
reg [32-1:0] arr_me3_f_global_v_wpv_e_0041=32'b11110100011011010111010001000000;
reg [32-1:0] arr_me3_f_global_v_wpv_e_0042=32'b11110100011110001010110101110101;
reg [32-1:0] arr_me3_f_global_v_wpv_e_0043=32'b11110100110000011100111000011111;
reg [32-1:0] arr_me3_f_global_v_wpv_e_0044=32'b11110100110001110001110011101101;
reg [32-1:0] arr_me3_f_global_v_wpv_e_0045=32'b11110100110011000011111111100000;
reg [32-1:0] arr_me3_f_global_v_wpv_e_0046=32'b11110100110100010011001111001101;
reg [32-1:0] arr_me3_f_global_v_wpv_e_0047=32'b11110100110101011111010110100101;
reg [32-1:0] arr_me3_f_global_v_wpv_e_0048=32'b11110100110110101000001001111010;
reg [32-1:0] arr_me3_f_global_v_wpv_e_0049=32'b11110100110111101101011101111101;
reg [32-1:0] arr_me3_f_global_v_wpv_e_0050=32'b11110100111000101111001000000010;
reg [32-1:0] arr_me3_f_global_v_wpv_e_0051=32'b11110100111001101100111110000001;
reg [32-1:0] arr_me3_f_global_v_wpv_e_0052=32'b11110100111010100110110110011001;
reg [32-1:0] arr_me3_f_global_v_wpv_e_0053=32'b11110100111011011100101000001101;
reg [32-1:0] arr_me3_f_global_v_wpv_e_0054=32'b11110100111100001110001011001100;
reg [32-1:0] arr_me3_f_global_v_wpv_e_0055=32'b11110100111100111011010111101100;
reg [32-1:0] arr_me3_f_global_v_wpv_e_0056=32'b11110100111101100100000110101111;
reg [32-1:0] arr_me3_f_global_v_wpv_e_0057=32'b11110100111110001000010010000100;
reg [32-1:0] arr_me3_f_global_v_wpv_e_0058=32'b11110100111110100111110100000110;
reg [32-1:0] arr_me3_f_global_v_wpv_e_0059=32'b11110100111111000010100111111100;
reg [32-1:0] arr_me3_f_global_v_wpv_e_0060=32'b11110100111111011000101001011111;
reg [32-1:0] arr_me3_f_global_v_wpv_e_0061=32'b11110100111111101001110101010110;
reg [32-1:0] arr_me3_f_global_v_wpv_e_0062=32'b11110100111111110110001000110111;
reg [32-1:0] arr_me3_f_global_v_wpv_e_0063=32'b11110100111111111101100010001000;
reg [32-1:0] arr_me3_f_global_v_wpv_i_e_0000=32'b01000000000000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_wpv_i_e_0001=32'b01110010111001000111110110011000;
reg [32-1:0] arr_me3_f_global_v_wpv_i_e_0002=32'b01110011011001000101111010011011;
reg [32-1:0] arr_me3_f_global_v_wpv_i_e_0003=32'b01110011110010110010000001000010;
reg [32-1:0] arr_me3_f_global_v_wpv_i_e_0004=32'b01110011111000111110001011100001;
reg [32-1:0] arr_me3_f_global_v_wpv_i_e_0005=32'b01110011111111000110011111100110;
reg [32-1:0] arr_me3_f_global_v_wpv_i_e_0006=32'b01110100010010100101000000011001;
reg [32-1:0] arr_me3_f_global_v_wpv_i_e_0007=32'b01110100010101100011111001101010;
reg [32-1:0] arr_me3_f_global_v_wpv_i_e_0008=32'b01110100011000011111011110001011;
reg [32-1:0] arr_me3_f_global_v_wpv_i_e_0009=32'b01110100011011010111010001000000;
reg [32-1:0] arr_me3_f_global_v_wpv_i_e_0010=32'b01110100011110001010110101110101;
reg [32-1:0] arr_me3_f_global_v_wpv_i_e_0011=32'b01110100110000011100111000011111;
reg [32-1:0] arr_me3_f_global_v_wpv_i_e_0012=32'b01110100110001110001110011101101;
reg [32-1:0] arr_me3_f_global_v_wpv_i_e_0013=32'b01110100110011000011111111100000;
reg [32-1:0] arr_me3_f_global_v_wpv_i_e_0014=32'b01110100110100010011001111001101;
reg [32-1:0] arr_me3_f_global_v_wpv_i_e_0015=32'b01110100110101011111010110100101;
reg [32-1:0] arr_me3_f_global_v_wpv_i_e_0016=32'b01110100110110101000001001111010;
reg [32-1:0] arr_me3_f_global_v_wpv_i_e_0017=32'b01110100110111101101011101111101;
reg [32-1:0] arr_me3_f_global_v_wpv_i_e_0018=32'b01110100111000101111001000000010;
reg [32-1:0] arr_me3_f_global_v_wpv_i_e_0019=32'b01110100111001101100111110000001;
reg [32-1:0] arr_me3_f_global_v_wpv_i_e_0020=32'b01110100111010100110110110011001;
reg [32-1:0] arr_me3_f_global_v_wpv_i_e_0021=32'b01110100111011011100101000001101;
reg [32-1:0] arr_me3_f_global_v_wpv_i_e_0022=32'b01110100111100001110001011001100;
reg [32-1:0] arr_me3_f_global_v_wpv_i_e_0023=32'b01110100111100111011010111101100;
reg [32-1:0] arr_me3_f_global_v_wpv_i_e_0024=32'b01110100111101100100000110101111;
reg [32-1:0] arr_me3_f_global_v_wpv_i_e_0025=32'b01110100111110001000010010000100;
reg [32-1:0] arr_me3_f_global_v_wpv_i_e_0026=32'b01110100111110100111110100000110;
reg [32-1:0] arr_me3_f_global_v_wpv_i_e_0027=32'b01110100111111000010100111111100;
reg [32-1:0] arr_me3_f_global_v_wpv_i_e_0028=32'b01110100111111011000101001011111;
reg [32-1:0] arr_me3_f_global_v_wpv_i_e_0029=32'b01110100111111101001110101010110;
reg [32-1:0] arr_me3_f_global_v_wpv_i_e_0030=32'b01110100111111110110001000110111;
reg [32-1:0] arr_me3_f_global_v_wpv_i_e_0031=32'b01110100111111111101100010001000;
reg [32-1:0] arr_me3_f_global_v_wpv_i_e_0032=32'b01110101010000000000000000000000;
reg [32-1:0] arr_me3_f_global_v_wpv_i_e_0033=32'b01110100111111111101100010001000;
reg [32-1:0] arr_me3_f_global_v_wpv_i_e_0034=32'b01110100111111110110001000110111;
reg [32-1:0] arr_me3_f_global_v_wpv_i_e_0035=32'b01110100111111101001110101010110;
reg [32-1:0] arr_me3_f_global_v_wpv_i_e_0036=32'b01110100111111011000101001011111;
reg [32-1:0] arr_me3_f_global_v_wpv_i_e_0037=32'b01110100111111000010100111111100;
reg [32-1:0] arr_me3_f_global_v_wpv_i_e_0038=32'b01110100111110100111110100000110;
reg [32-1:0] arr_me3_f_global_v_wpv_i_e_0039=32'b01110100111110001000010010000100;
reg [32-1:0] arr_me3_f_global_v_wpv_i_e_0040=32'b01110100111101100100000110101111;
reg [32-1:0] arr_me3_f_global_v_wpv_i_e_0041=32'b01110100111100111011010111101100;
reg [32-1:0] arr_me3_f_global_v_wpv_i_e_0042=32'b01110100111100001110001011001100;
reg [32-1:0] arr_me3_f_global_v_wpv_i_e_0043=32'b01110100111011011100101000001101;
reg [32-1:0] arr_me3_f_global_v_wpv_i_e_0044=32'b01110100111010100110110110011001;
reg [32-1:0] arr_me3_f_global_v_wpv_i_e_0045=32'b01110100111001101100111110000001;
reg [32-1:0] arr_me3_f_global_v_wpv_i_e_0046=32'b01110100111000101111001000000010;
reg [32-1:0] arr_me3_f_global_v_wpv_i_e_0047=32'b01110100110111101101011101111101;
reg [32-1:0] arr_me3_f_global_v_wpv_i_e_0048=32'b01110100110110101000001001111010;
reg [32-1:0] arr_me3_f_global_v_wpv_i_e_0049=32'b01110100110101011111010110100101;
reg [32-1:0] arr_me3_f_global_v_wpv_i_e_0050=32'b01110100110100010011001111001101;
reg [32-1:0] arr_me3_f_global_v_wpv_i_e_0051=32'b01110100110011000011111111100000;
reg [32-1:0] arr_me3_f_global_v_wpv_i_e_0052=32'b01110100110001110001110011101101;
reg [32-1:0] arr_me3_f_global_v_wpv_i_e_0053=32'b01110100110000011100111000011111;
reg [32-1:0] arr_me3_f_global_v_wpv_i_e_0054=32'b01110100011110001010110101110101;
reg [32-1:0] arr_me3_f_global_v_wpv_i_e_0055=32'b01110100011011010111010001000000;
reg [32-1:0] arr_me3_f_global_v_wpv_i_e_0056=32'b01110100011000011111011110001011;
reg [32-1:0] arr_me3_f_global_v_wpv_i_e_0057=32'b01110100010101100011111001101010;
reg [32-1:0] arr_me3_f_global_v_wpv_i_e_0058=32'b01110100010010100101000000011001;
reg [32-1:0] arr_me3_f_global_v_wpv_i_e_0059=32'b01110011111111000110011111100110;
reg [32-1:0] arr_me3_f_global_v_wpv_i_e_0060=32'b01110011111000111110001011100001;
reg [32-1:0] arr_me3_f_global_v_wpv_i_e_0061=32'b01110011110010110010000001000010;
reg [32-1:0] arr_me3_f_global_v_wpv_i_e_0062=32'b01110011011001000101111010011011;
reg [32-1:0] arr_me3_f_global_v_wpv_i_e_0063=32'b01110010111001000111110110011000;
integer sm_me2; always @ (*) sm_me2 = (out[31]) ? -out[22:0] : out[22:0];
integer  e_me2; always @ (*)  e_me2 = $signed(out[30:23]);
real arr_me2_f_main_v_output_buffer_real_e_0000 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0001 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0002 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0003 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0004 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0005 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0006 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0007 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0008 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0009 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0010 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0011 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0012 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0013 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0014 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0015 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0016 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0017 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0018 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0019 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0020 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0021 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0022 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0023 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0024 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0025 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0026 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0027 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0028 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0029 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0030 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0031 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0032 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0033 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0034 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0035 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0036 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0037 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0038 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0039 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0040 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0041 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0042 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0043 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0044 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0045 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0046 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0047 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0048 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0049 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0050 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0051 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0052 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0053 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0054 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0055 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0056 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0057 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0058 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0059 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0060 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0061 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0062 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0063 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0064 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0065 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0066 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0067 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0068 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0069 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0070 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0071 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0072 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0073 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0074 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0075 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0076 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0077 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0078 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0079 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0080 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0081 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0082 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0083 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0084 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0085 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0086 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0087 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0088 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0089 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0090 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0091 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0092 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0093 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0094 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0095 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0096 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0097 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0098 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0099 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0100 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0101 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0102 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0103 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0104 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0105 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0106 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0107 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0108 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0109 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0110 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0111 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0112 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0113 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0114 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0115 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0116 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0117 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0118 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0119 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0120 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0121 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0122 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0123 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0124 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0125 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0126 = 0.000000;
real arr_me2_f_main_v_output_buffer_real_e_0127 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0000 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0001 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0002 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0003 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0004 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0005 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0006 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0007 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0008 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0009 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0010 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0011 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0012 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0013 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0014 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0015 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0016 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0017 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0018 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0019 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0020 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0021 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0022 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0023 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0024 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0025 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0026 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0027 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0028 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0029 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0030 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0031 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0032 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0033 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0034 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0035 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0036 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0037 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0038 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0039 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0040 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0041 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0042 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0043 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0044 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0045 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0046 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0047 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0048 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0049 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0050 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0051 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0052 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0053 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0054 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0055 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0056 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0057 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0058 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0059 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0060 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0061 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0062 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0063 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0064 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0065 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0066 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0067 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0068 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0069 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0070 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0071 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0072 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0073 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0074 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0075 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0076 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0077 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0078 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0079 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0080 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0081 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0082 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0083 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0084 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0085 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0086 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0087 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0088 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0089 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0090 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0091 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0092 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0093 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0094 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0095 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0096 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0097 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0098 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0099 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0100 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0101 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0102 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0103 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0104 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0105 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0106 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0107 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0108 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0109 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0110 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0111 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0112 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0113 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0114 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0115 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0116 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0117 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0118 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0119 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0120 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0121 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0122 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0123 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0124 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0125 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0126 = 0.000000;
real arr_me2_f_main_v_output_buffer_imag_e_0127 = 0.000000;
real arr_me2_f_main_v_buffer_e_0000 = 0.000000;
real arr_me2_f_main_v_buffer_e_0001 = 0.000000;
real arr_me2_f_main_v_buffer_e_0002 = 0.000000;
real arr_me2_f_main_v_buffer_e_0003 = 0.000000;
real arr_me2_f_main_v_buffer_e_0004 = 0.000000;
real arr_me2_f_main_v_buffer_e_0005 = 0.000000;
real arr_me2_f_main_v_buffer_e_0006 = 0.000000;
real arr_me2_f_main_v_buffer_e_0007 = 0.000000;
real arr_me2_f_main_v_buffer_e_0008 = 0.000000;
real arr_me2_f_main_v_buffer_e_0009 = 0.000000;
real arr_me2_f_main_v_buffer_e_0010 = 0.000000;
real arr_me2_f_main_v_buffer_e_0011 = 0.000000;
real arr_me2_f_main_v_buffer_e_0012 = 0.000000;
real arr_me2_f_main_v_buffer_e_0013 = 0.000000;
real arr_me2_f_main_v_buffer_e_0014 = 0.000000;
real arr_me2_f_main_v_buffer_e_0015 = 0.000000;
real arr_me2_f_main_v_buffer_e_0016 = 0.000000;
real arr_me2_f_main_v_buffer_e_0017 = 0.000000;
real arr_me2_f_main_v_buffer_e_0018 = 0.000000;
real arr_me2_f_main_v_buffer_e_0019 = 0.000000;
real arr_me2_f_main_v_buffer_e_0020 = 0.000000;
real arr_me2_f_main_v_buffer_e_0021 = 0.000000;
real arr_me2_f_main_v_buffer_e_0022 = 0.000000;
real arr_me2_f_main_v_buffer_e_0023 = 0.000000;
real arr_me2_f_main_v_buffer_e_0024 = 0.000000;
real arr_me2_f_main_v_buffer_e_0025 = 0.000000;
real arr_me2_f_main_v_buffer_e_0026 = 0.000000;
real arr_me2_f_main_v_buffer_e_0027 = 0.000000;
real arr_me2_f_main_v_buffer_e_0028 = 0.000000;
real arr_me2_f_main_v_buffer_e_0029 = 0.000000;
real arr_me2_f_main_v_buffer_e_0030 = 0.000000;
real arr_me2_f_main_v_buffer_e_0031 = 0.000000;
real arr_me2_f_main_v_buffer_e_0032 = 0.000000;
real arr_me2_f_main_v_buffer_e_0033 = 0.000000;
real arr_me2_f_main_v_buffer_e_0034 = 0.000000;
real arr_me2_f_main_v_buffer_e_0035 = 0.000000;
real arr_me2_f_main_v_buffer_e_0036 = 0.000000;
real arr_me2_f_main_v_buffer_e_0037 = 0.000000;
real arr_me2_f_main_v_buffer_e_0038 = 0.000000;
real arr_me2_f_main_v_buffer_e_0039 = 0.000000;
real arr_me2_f_main_v_buffer_e_0040 = 0.000000;
real arr_me2_f_main_v_buffer_e_0041 = 0.000000;
real arr_me2_f_main_v_buffer_e_0042 = 0.000000;
real arr_me2_f_main_v_buffer_e_0043 = 0.000000;
real arr_me2_f_main_v_buffer_e_0044 = 0.000000;
real arr_me2_f_main_v_buffer_e_0045 = 0.000000;
real arr_me2_f_main_v_buffer_e_0046 = 0.000000;
real arr_me2_f_main_v_buffer_e_0047 = 0.000000;
real arr_me2_f_main_v_buffer_e_0048 = 0.000000;
real arr_me2_f_main_v_buffer_e_0049 = 0.000000;
real arr_me2_f_main_v_buffer_e_0050 = 0.000000;
real arr_me2_f_main_v_buffer_e_0051 = 0.000000;
real arr_me2_f_main_v_buffer_e_0052 = 0.000000;
real arr_me2_f_main_v_buffer_e_0053 = 0.000000;
real arr_me2_f_main_v_buffer_e_0054 = 0.000000;
real arr_me2_f_main_v_buffer_e_0055 = 0.000000;
real arr_me2_f_main_v_buffer_e_0056 = 0.000000;
real arr_me2_f_main_v_buffer_e_0057 = 0.000000;
real arr_me2_f_main_v_buffer_e_0058 = 0.000000;
real arr_me2_f_main_v_buffer_e_0059 = 0.000000;
real arr_me2_f_main_v_buffer_e_0060 = 0.000000;
real arr_me2_f_main_v_buffer_e_0061 = 0.000000;
real arr_me2_f_main_v_buffer_e_0062 = 0.000000;
real arr_me2_f_main_v_buffer_e_0063 = 0.000000;
real arr_me2_f_main_v_buffer_e_0064 = 0.000000;
real arr_me2_f_main_v_buffer_e_0065 = 0.000000;
real arr_me2_f_main_v_buffer_e_0066 = 0.000000;
real arr_me2_f_main_v_buffer_e_0067 = 0.000000;
real arr_me2_f_main_v_buffer_e_0068 = 0.000000;
real arr_me2_f_main_v_buffer_e_0069 = 0.000000;
real arr_me2_f_main_v_buffer_e_0070 = 0.000000;
real arr_me2_f_main_v_buffer_e_0071 = 0.000000;
real arr_me2_f_main_v_buffer_e_0072 = 0.000000;
real arr_me2_f_main_v_buffer_e_0073 = 0.000000;
real arr_me2_f_main_v_buffer_e_0074 = 0.000000;
real arr_me2_f_main_v_buffer_e_0075 = 0.000000;
real arr_me2_f_main_v_buffer_e_0076 = 0.000000;
real arr_me2_f_main_v_buffer_e_0077 = 0.000000;
real arr_me2_f_main_v_buffer_e_0078 = 0.000000;
real arr_me2_f_main_v_buffer_e_0079 = 0.000000;
real arr_me2_f_main_v_buffer_e_0080 = 0.000000;
real arr_me2_f_main_v_buffer_e_0081 = 0.000000;
real arr_me2_f_main_v_buffer_e_0082 = 0.000000;
real arr_me2_f_main_v_buffer_e_0083 = 0.000000;
real arr_me2_f_main_v_buffer_e_0084 = 0.000000;
real arr_me2_f_main_v_buffer_e_0085 = 0.000000;
real arr_me2_f_main_v_buffer_e_0086 = 0.000000;
real arr_me2_f_main_v_buffer_e_0087 = 0.000000;
real arr_me2_f_main_v_buffer_e_0088 = 0.000000;
real arr_me2_f_main_v_buffer_e_0089 = 0.000000;
real arr_me2_f_main_v_buffer_e_0090 = 0.000000;
real arr_me2_f_main_v_buffer_e_0091 = 0.000000;
real arr_me2_f_main_v_buffer_e_0092 = 0.000000;
real arr_me2_f_main_v_buffer_e_0093 = 0.000000;
real arr_me2_f_main_v_buffer_e_0094 = 0.000000;
real arr_me2_f_main_v_buffer_e_0095 = 0.000000;
real arr_me2_f_main_v_buffer_e_0096 = 0.000000;
real arr_me2_f_main_v_buffer_e_0097 = 0.000000;
real arr_me2_f_main_v_buffer_e_0098 = 0.000000;
real arr_me2_f_main_v_buffer_e_0099 = 0.000000;
real arr_me2_f_main_v_buffer_e_0100 = 0.000000;
real arr_me2_f_main_v_buffer_e_0101 = 0.000000;
real arr_me2_f_main_v_buffer_e_0102 = 0.000000;
real arr_me2_f_main_v_buffer_e_0103 = 0.000000;
real arr_me2_f_main_v_buffer_e_0104 = 0.000000;
real arr_me2_f_main_v_buffer_e_0105 = 0.000000;
real arr_me2_f_main_v_buffer_e_0106 = 0.000000;
real arr_me2_f_main_v_buffer_e_0107 = 0.000000;
real arr_me2_f_main_v_buffer_e_0108 = 0.000000;
real arr_me2_f_main_v_buffer_e_0109 = 0.000000;
real arr_me2_f_main_v_buffer_e_0110 = 0.000000;
real arr_me2_f_main_v_buffer_e_0111 = 0.000000;
real arr_me2_f_main_v_buffer_e_0112 = 0.000000;
real arr_me2_f_main_v_buffer_e_0113 = 0.000000;
real arr_me2_f_main_v_buffer_e_0114 = 0.000000;
real arr_me2_f_main_v_buffer_e_0115 = 0.000000;
real arr_me2_f_main_v_buffer_e_0116 = 0.000000;
real arr_me2_f_main_v_buffer_e_0117 = 0.000000;
real arr_me2_f_main_v_buffer_e_0118 = 0.000000;
real arr_me2_f_main_v_buffer_e_0119 = 0.000000;
real arr_me2_f_main_v_buffer_e_0120 = 0.000000;
real arr_me2_f_main_v_buffer_e_0121 = 0.000000;
real arr_me2_f_main_v_buffer_e_0122 = 0.000000;
real arr_me2_f_main_v_buffer_e_0123 = 0.000000;
real arr_me2_f_main_v_buffer_e_0124 = 0.000000;
real arr_me2_f_main_v_buffer_e_0125 = 0.000000;
real arr_me2_f_main_v_buffer_e_0126 = 0.000000;
real arr_me2_f_main_v_buffer_e_0127 = 0.000000;

always @ (posedge clk) begin
   if (mem_addr_wr == 0 && mem_wr) arr_me3_f_global_v_E0_e_0000 <= out;
   if (mem_addr_wr == 1 && mem_wr) arr_me3_f_global_v_E0_e_0001 <= out;
   if (mem_addr_wr == 2 && mem_wr) arr_me3_f_global_v_E0_e_0002 <= out;
   if (mem_addr_wr == 3 && mem_wr) arr_me3_f_global_v_E0_e_0003 <= out;
   if (mem_addr_wr == 4 && mem_wr) arr_me3_f_global_v_E0_e_0004 <= out;
   if (mem_addr_wr == 5 && mem_wr) arr_me3_f_global_v_E0_e_0005 <= out;
   if (mem_addr_wr == 6 && mem_wr) arr_me3_f_global_v_E0_e_0006 <= out;
   if (mem_addr_wr == 7 && mem_wr) arr_me3_f_global_v_E0_e_0007 <= out;
   if (mem_addr_wr == 8 && mem_wr) arr_me3_f_global_v_E0_e_0008 <= out;
   if (mem_addr_wr == 9 && mem_wr) arr_me3_f_global_v_E0_e_0009 <= out;
   if (mem_addr_wr == 10 && mem_wr) arr_me3_f_global_v_E0_e_0010 <= out;
   if (mem_addr_wr == 11 && mem_wr) arr_me3_f_global_v_E0_e_0011 <= out;
   if (mem_addr_wr == 12 && mem_wr) arr_me3_f_global_v_E0_e_0012 <= out;
   if (mem_addr_wr == 13 && mem_wr) arr_me3_f_global_v_E0_e_0013 <= out;
   if (mem_addr_wr == 14 && mem_wr) arr_me3_f_global_v_E0_e_0014 <= out;
   if (mem_addr_wr == 15 && mem_wr) arr_me3_f_global_v_E0_e_0015 <= out;
   if (mem_addr_wr == 16 && mem_wr) arr_me3_f_global_v_E0_e_0016 <= out;
   if (mem_addr_wr == 17 && mem_wr) arr_me3_f_global_v_E0_e_0017 <= out;
   if (mem_addr_wr == 18 && mem_wr) arr_me3_f_global_v_E0_e_0018 <= out;
   if (mem_addr_wr == 19 && mem_wr) arr_me3_f_global_v_E0_e_0019 <= out;
   if (mem_addr_wr == 20 && mem_wr) arr_me3_f_global_v_E0_e_0020 <= out;
   if (mem_addr_wr == 21 && mem_wr) arr_me3_f_global_v_E0_e_0021 <= out;
   if (mem_addr_wr == 22 && mem_wr) arr_me3_f_global_v_E0_e_0022 <= out;
   if (mem_addr_wr == 23 && mem_wr) arr_me3_f_global_v_E0_e_0023 <= out;
   if (mem_addr_wr == 24 && mem_wr) arr_me3_f_global_v_E0_e_0024 <= out;
   if (mem_addr_wr == 25 && mem_wr) arr_me3_f_global_v_E0_e_0025 <= out;
   if (mem_addr_wr == 26 && mem_wr) arr_me3_f_global_v_E0_e_0026 <= out;
   if (mem_addr_wr == 27 && mem_wr) arr_me3_f_global_v_E0_e_0027 <= out;
   if (mem_addr_wr == 28 && mem_wr) arr_me3_f_global_v_E0_e_0028 <= out;
   if (mem_addr_wr == 29 && mem_wr) arr_me3_f_global_v_E0_e_0029 <= out;
   if (mem_addr_wr == 30 && mem_wr) arr_me3_f_global_v_E0_e_0030 <= out;
   if (mem_addr_wr == 31 && mem_wr) arr_me3_f_global_v_E0_e_0031 <= out;
   if (mem_addr_wr == 32 && mem_wr) arr_me3_f_global_v_E0_e_0032 <= out;
   if (mem_addr_wr == 33 && mem_wr) arr_me3_f_global_v_E0_e_0033 <= out;
   if (mem_addr_wr == 34 && mem_wr) arr_me3_f_global_v_E0_e_0034 <= out;
   if (mem_addr_wr == 35 && mem_wr) arr_me3_f_global_v_E0_e_0035 <= out;
   if (mem_addr_wr == 36 && mem_wr) arr_me3_f_global_v_E0_e_0036 <= out;
   if (mem_addr_wr == 37 && mem_wr) arr_me3_f_global_v_E0_e_0037 <= out;
   if (mem_addr_wr == 38 && mem_wr) arr_me3_f_global_v_E0_e_0038 <= out;
   if (mem_addr_wr == 39 && mem_wr) arr_me3_f_global_v_E0_e_0039 <= out;
   if (mem_addr_wr == 40 && mem_wr) arr_me3_f_global_v_E0_e_0040 <= out;
   if (mem_addr_wr == 41 && mem_wr) arr_me3_f_global_v_E0_e_0041 <= out;
   if (mem_addr_wr == 42 && mem_wr) arr_me3_f_global_v_E0_e_0042 <= out;
   if (mem_addr_wr == 43 && mem_wr) arr_me3_f_global_v_E0_e_0043 <= out;
   if (mem_addr_wr == 44 && mem_wr) arr_me3_f_global_v_E0_e_0044 <= out;
   if (mem_addr_wr == 45 && mem_wr) arr_me3_f_global_v_E0_e_0045 <= out;
   if (mem_addr_wr == 46 && mem_wr) arr_me3_f_global_v_E0_e_0046 <= out;
   if (mem_addr_wr == 47 && mem_wr) arr_me3_f_global_v_E0_e_0047 <= out;
   if (mem_addr_wr == 48 && mem_wr) arr_me3_f_global_v_E0_e_0048 <= out;
   if (mem_addr_wr == 49 && mem_wr) arr_me3_f_global_v_E0_e_0049 <= out;
   if (mem_addr_wr == 50 && mem_wr) arr_me3_f_global_v_E0_e_0050 <= out;
   if (mem_addr_wr == 51 && mem_wr) arr_me3_f_global_v_E0_e_0051 <= out;
   if (mem_addr_wr == 52 && mem_wr) arr_me3_f_global_v_E0_e_0052 <= out;
   if (mem_addr_wr == 53 && mem_wr) arr_me3_f_global_v_E0_e_0053 <= out;
   if (mem_addr_wr == 54 && mem_wr) arr_me3_f_global_v_E0_e_0054 <= out;
   if (mem_addr_wr == 55 && mem_wr) arr_me3_f_global_v_E0_e_0055 <= out;
   if (mem_addr_wr == 56 && mem_wr) arr_me3_f_global_v_E0_e_0056 <= out;
   if (mem_addr_wr == 57 && mem_wr) arr_me3_f_global_v_E0_e_0057 <= out;
   if (mem_addr_wr == 58 && mem_wr) arr_me3_f_global_v_E0_e_0058 <= out;
   if (mem_addr_wr == 59 && mem_wr) arr_me3_f_global_v_E0_e_0059 <= out;
   if (mem_addr_wr == 60 && mem_wr) arr_me3_f_global_v_E0_e_0060 <= out;
   if (mem_addr_wr == 61 && mem_wr) arr_me3_f_global_v_E0_e_0061 <= out;
   if (mem_addr_wr == 62 && mem_wr) arr_me3_f_global_v_E0_e_0062 <= out;
   if (mem_addr_wr == 63 && mem_wr) arr_me3_f_global_v_E0_e_0063 <= out;
   if (mem_addr_wr == 64 && mem_wr) arr_me3_f_global_v_E0_e_0064 <= out;
   if (mem_addr_wr == 65 && mem_wr) arr_me3_f_global_v_E0_e_0065 <= out;
   if (mem_addr_wr == 66 && mem_wr) arr_me3_f_global_v_E0_e_0066 <= out;
   if (mem_addr_wr == 67 && mem_wr) arr_me3_f_global_v_E0_e_0067 <= out;
   if (mem_addr_wr == 68 && mem_wr) arr_me3_f_global_v_E0_e_0068 <= out;
   if (mem_addr_wr == 69 && mem_wr) arr_me3_f_global_v_E0_e_0069 <= out;
   if (mem_addr_wr == 70 && mem_wr) arr_me3_f_global_v_E0_e_0070 <= out;
   if (mem_addr_wr == 71 && mem_wr) arr_me3_f_global_v_E0_e_0071 <= out;
   if (mem_addr_wr == 72 && mem_wr) arr_me3_f_global_v_E0_e_0072 <= out;
   if (mem_addr_wr == 73 && mem_wr) arr_me3_f_global_v_E0_e_0073 <= out;
   if (mem_addr_wr == 74 && mem_wr) arr_me3_f_global_v_E0_e_0074 <= out;
   if (mem_addr_wr == 75 && mem_wr) arr_me3_f_global_v_E0_e_0075 <= out;
   if (mem_addr_wr == 76 && mem_wr) arr_me3_f_global_v_E0_e_0076 <= out;
   if (mem_addr_wr == 77 && mem_wr) arr_me3_f_global_v_E0_e_0077 <= out;
   if (mem_addr_wr == 78 && mem_wr) arr_me3_f_global_v_E0_e_0078 <= out;
   if (mem_addr_wr == 79 && mem_wr) arr_me3_f_global_v_E0_e_0079 <= out;
   if (mem_addr_wr == 80 && mem_wr) arr_me3_f_global_v_E0_e_0080 <= out;
   if (mem_addr_wr == 81 && mem_wr) arr_me3_f_global_v_E0_e_0081 <= out;
   if (mem_addr_wr == 82 && mem_wr) arr_me3_f_global_v_E0_e_0082 <= out;
   if (mem_addr_wr == 83 && mem_wr) arr_me3_f_global_v_E0_e_0083 <= out;
   if (mem_addr_wr == 84 && mem_wr) arr_me3_f_global_v_E0_e_0084 <= out;
   if (mem_addr_wr == 85 && mem_wr) arr_me3_f_global_v_E0_e_0085 <= out;
   if (mem_addr_wr == 86 && mem_wr) arr_me3_f_global_v_E0_e_0086 <= out;
   if (mem_addr_wr == 87 && mem_wr) arr_me3_f_global_v_E0_e_0087 <= out;
   if (mem_addr_wr == 88 && mem_wr) arr_me3_f_global_v_E0_e_0088 <= out;
   if (mem_addr_wr == 89 && mem_wr) arr_me3_f_global_v_E0_e_0089 <= out;
   if (mem_addr_wr == 90 && mem_wr) arr_me3_f_global_v_E0_e_0090 <= out;
   if (mem_addr_wr == 91 && mem_wr) arr_me3_f_global_v_E0_e_0091 <= out;
   if (mem_addr_wr == 92 && mem_wr) arr_me3_f_global_v_E0_e_0092 <= out;
   if (mem_addr_wr == 93 && mem_wr) arr_me3_f_global_v_E0_e_0093 <= out;
   if (mem_addr_wr == 94 && mem_wr) arr_me3_f_global_v_E0_e_0094 <= out;
   if (mem_addr_wr == 95 && mem_wr) arr_me3_f_global_v_E0_e_0095 <= out;
   if (mem_addr_wr == 96 && mem_wr) arr_me3_f_global_v_E0_e_0096 <= out;
   if (mem_addr_wr == 97 && mem_wr) arr_me3_f_global_v_E0_e_0097 <= out;
   if (mem_addr_wr == 98 && mem_wr) arr_me3_f_global_v_E0_e_0098 <= out;
   if (mem_addr_wr == 99 && mem_wr) arr_me3_f_global_v_E0_e_0099 <= out;
   if (mem_addr_wr == 100 && mem_wr) arr_me3_f_global_v_E0_e_0100 <= out;
   if (mem_addr_wr == 101 && mem_wr) arr_me3_f_global_v_E0_e_0101 <= out;
   if (mem_addr_wr == 102 && mem_wr) arr_me3_f_global_v_E0_e_0102 <= out;
   if (mem_addr_wr == 103 && mem_wr) arr_me3_f_global_v_E0_e_0103 <= out;
   if (mem_addr_wr == 104 && mem_wr) arr_me3_f_global_v_E0_e_0104 <= out;
   if (mem_addr_wr == 105 && mem_wr) arr_me3_f_global_v_E0_e_0105 <= out;
   if (mem_addr_wr == 106 && mem_wr) arr_me3_f_global_v_E0_e_0106 <= out;
   if (mem_addr_wr == 107 && mem_wr) arr_me3_f_global_v_E0_e_0107 <= out;
   if (mem_addr_wr == 108 && mem_wr) arr_me3_f_global_v_E0_e_0108 <= out;
   if (mem_addr_wr == 109 && mem_wr) arr_me3_f_global_v_E0_e_0109 <= out;
   if (mem_addr_wr == 110 && mem_wr) arr_me3_f_global_v_E0_e_0110 <= out;
   if (mem_addr_wr == 111 && mem_wr) arr_me3_f_global_v_E0_e_0111 <= out;
   if (mem_addr_wr == 112 && mem_wr) arr_me3_f_global_v_E0_e_0112 <= out;
   if (mem_addr_wr == 113 && mem_wr) arr_me3_f_global_v_E0_e_0113 <= out;
   if (mem_addr_wr == 114 && mem_wr) arr_me3_f_global_v_E0_e_0114 <= out;
   if (mem_addr_wr == 115 && mem_wr) arr_me3_f_global_v_E0_e_0115 <= out;
   if (mem_addr_wr == 116 && mem_wr) arr_me3_f_global_v_E0_e_0116 <= out;
   if (mem_addr_wr == 117 && mem_wr) arr_me3_f_global_v_E0_e_0117 <= out;
   if (mem_addr_wr == 118 && mem_wr) arr_me3_f_global_v_E0_e_0118 <= out;
   if (mem_addr_wr == 119 && mem_wr) arr_me3_f_global_v_E0_e_0119 <= out;
   if (mem_addr_wr == 120 && mem_wr) arr_me3_f_global_v_E0_e_0120 <= out;
   if (mem_addr_wr == 121 && mem_wr) arr_me3_f_global_v_E0_e_0121 <= out;
   if (mem_addr_wr == 122 && mem_wr) arr_me3_f_global_v_E0_e_0122 <= out;
   if (mem_addr_wr == 123 && mem_wr) arr_me3_f_global_v_E0_e_0123 <= out;
   if (mem_addr_wr == 124 && mem_wr) arr_me3_f_global_v_E0_e_0124 <= out;
   if (mem_addr_wr == 125 && mem_wr) arr_me3_f_global_v_E0_e_0125 <= out;
   if (mem_addr_wr == 126 && mem_wr) arr_me3_f_global_v_E0_e_0126 <= out;
   if (mem_addr_wr == 127 && mem_wr) arr_me3_f_global_v_E0_e_0127 <= out;
   if (mem_addr_wr == 128 && mem_wr) arr_me3_f_global_v_E0_i_e_0000 <= out;
   if (mem_addr_wr == 129 && mem_wr) arr_me3_f_global_v_E0_i_e_0001 <= out;
   if (mem_addr_wr == 130 && mem_wr) arr_me3_f_global_v_E0_i_e_0002 <= out;
   if (mem_addr_wr == 131 && mem_wr) arr_me3_f_global_v_E0_i_e_0003 <= out;
   if (mem_addr_wr == 132 && mem_wr) arr_me3_f_global_v_E0_i_e_0004 <= out;
   if (mem_addr_wr == 133 && mem_wr) arr_me3_f_global_v_E0_i_e_0005 <= out;
   if (mem_addr_wr == 134 && mem_wr) arr_me3_f_global_v_E0_i_e_0006 <= out;
   if (mem_addr_wr == 135 && mem_wr) arr_me3_f_global_v_E0_i_e_0007 <= out;
   if (mem_addr_wr == 136 && mem_wr) arr_me3_f_global_v_E0_i_e_0008 <= out;
   if (mem_addr_wr == 137 && mem_wr) arr_me3_f_global_v_E0_i_e_0009 <= out;
   if (mem_addr_wr == 138 && mem_wr) arr_me3_f_global_v_E0_i_e_0010 <= out;
   if (mem_addr_wr == 139 && mem_wr) arr_me3_f_global_v_E0_i_e_0011 <= out;
   if (mem_addr_wr == 140 && mem_wr) arr_me3_f_global_v_E0_i_e_0012 <= out;
   if (mem_addr_wr == 141 && mem_wr) arr_me3_f_global_v_E0_i_e_0013 <= out;
   if (mem_addr_wr == 142 && mem_wr) arr_me3_f_global_v_E0_i_e_0014 <= out;
   if (mem_addr_wr == 143 && mem_wr) arr_me3_f_global_v_E0_i_e_0015 <= out;
   if (mem_addr_wr == 144 && mem_wr) arr_me3_f_global_v_E0_i_e_0016 <= out;
   if (mem_addr_wr == 145 && mem_wr) arr_me3_f_global_v_E0_i_e_0017 <= out;
   if (mem_addr_wr == 146 && mem_wr) arr_me3_f_global_v_E0_i_e_0018 <= out;
   if (mem_addr_wr == 147 && mem_wr) arr_me3_f_global_v_E0_i_e_0019 <= out;
   if (mem_addr_wr == 148 && mem_wr) arr_me3_f_global_v_E0_i_e_0020 <= out;
   if (mem_addr_wr == 149 && mem_wr) arr_me3_f_global_v_E0_i_e_0021 <= out;
   if (mem_addr_wr == 150 && mem_wr) arr_me3_f_global_v_E0_i_e_0022 <= out;
   if (mem_addr_wr == 151 && mem_wr) arr_me3_f_global_v_E0_i_e_0023 <= out;
   if (mem_addr_wr == 152 && mem_wr) arr_me3_f_global_v_E0_i_e_0024 <= out;
   if (mem_addr_wr == 153 && mem_wr) arr_me3_f_global_v_E0_i_e_0025 <= out;
   if (mem_addr_wr == 154 && mem_wr) arr_me3_f_global_v_E0_i_e_0026 <= out;
   if (mem_addr_wr == 155 && mem_wr) arr_me3_f_global_v_E0_i_e_0027 <= out;
   if (mem_addr_wr == 156 && mem_wr) arr_me3_f_global_v_E0_i_e_0028 <= out;
   if (mem_addr_wr == 157 && mem_wr) arr_me3_f_global_v_E0_i_e_0029 <= out;
   if (mem_addr_wr == 158 && mem_wr) arr_me3_f_global_v_E0_i_e_0030 <= out;
   if (mem_addr_wr == 159 && mem_wr) arr_me3_f_global_v_E0_i_e_0031 <= out;
   if (mem_addr_wr == 160 && mem_wr) arr_me3_f_global_v_E0_i_e_0032 <= out;
   if (mem_addr_wr == 161 && mem_wr) arr_me3_f_global_v_E0_i_e_0033 <= out;
   if (mem_addr_wr == 162 && mem_wr) arr_me3_f_global_v_E0_i_e_0034 <= out;
   if (mem_addr_wr == 163 && mem_wr) arr_me3_f_global_v_E0_i_e_0035 <= out;
   if (mem_addr_wr == 164 && mem_wr) arr_me3_f_global_v_E0_i_e_0036 <= out;
   if (mem_addr_wr == 165 && mem_wr) arr_me3_f_global_v_E0_i_e_0037 <= out;
   if (mem_addr_wr == 166 && mem_wr) arr_me3_f_global_v_E0_i_e_0038 <= out;
   if (mem_addr_wr == 167 && mem_wr) arr_me3_f_global_v_E0_i_e_0039 <= out;
   if (mem_addr_wr == 168 && mem_wr) arr_me3_f_global_v_E0_i_e_0040 <= out;
   if (mem_addr_wr == 169 && mem_wr) arr_me3_f_global_v_E0_i_e_0041 <= out;
   if (mem_addr_wr == 170 && mem_wr) arr_me3_f_global_v_E0_i_e_0042 <= out;
   if (mem_addr_wr == 171 && mem_wr) arr_me3_f_global_v_E0_i_e_0043 <= out;
   if (mem_addr_wr == 172 && mem_wr) arr_me3_f_global_v_E0_i_e_0044 <= out;
   if (mem_addr_wr == 173 && mem_wr) arr_me3_f_global_v_E0_i_e_0045 <= out;
   if (mem_addr_wr == 174 && mem_wr) arr_me3_f_global_v_E0_i_e_0046 <= out;
   if (mem_addr_wr == 175 && mem_wr) arr_me3_f_global_v_E0_i_e_0047 <= out;
   if (mem_addr_wr == 176 && mem_wr) arr_me3_f_global_v_E0_i_e_0048 <= out;
   if (mem_addr_wr == 177 && mem_wr) arr_me3_f_global_v_E0_i_e_0049 <= out;
   if (mem_addr_wr == 178 && mem_wr) arr_me3_f_global_v_E0_i_e_0050 <= out;
   if (mem_addr_wr == 179 && mem_wr) arr_me3_f_global_v_E0_i_e_0051 <= out;
   if (mem_addr_wr == 180 && mem_wr) arr_me3_f_global_v_E0_i_e_0052 <= out;
   if (mem_addr_wr == 181 && mem_wr) arr_me3_f_global_v_E0_i_e_0053 <= out;
   if (mem_addr_wr == 182 && mem_wr) arr_me3_f_global_v_E0_i_e_0054 <= out;
   if (mem_addr_wr == 183 && mem_wr) arr_me3_f_global_v_E0_i_e_0055 <= out;
   if (mem_addr_wr == 184 && mem_wr) arr_me3_f_global_v_E0_i_e_0056 <= out;
   if (mem_addr_wr == 185 && mem_wr) arr_me3_f_global_v_E0_i_e_0057 <= out;
   if (mem_addr_wr == 186 && mem_wr) arr_me3_f_global_v_E0_i_e_0058 <= out;
   if (mem_addr_wr == 187 && mem_wr) arr_me3_f_global_v_E0_i_e_0059 <= out;
   if (mem_addr_wr == 188 && mem_wr) arr_me3_f_global_v_E0_i_e_0060 <= out;
   if (mem_addr_wr == 189 && mem_wr) arr_me3_f_global_v_E0_i_e_0061 <= out;
   if (mem_addr_wr == 190 && mem_wr) arr_me3_f_global_v_E0_i_e_0062 <= out;
   if (mem_addr_wr == 191 && mem_wr) arr_me3_f_global_v_E0_i_e_0063 <= out;
   if (mem_addr_wr == 192 && mem_wr) arr_me3_f_global_v_E0_i_e_0064 <= out;
   if (mem_addr_wr == 193 && mem_wr) arr_me3_f_global_v_E0_i_e_0065 <= out;
   if (mem_addr_wr == 194 && mem_wr) arr_me3_f_global_v_E0_i_e_0066 <= out;
   if (mem_addr_wr == 195 && mem_wr) arr_me3_f_global_v_E0_i_e_0067 <= out;
   if (mem_addr_wr == 196 && mem_wr) arr_me3_f_global_v_E0_i_e_0068 <= out;
   if (mem_addr_wr == 197 && mem_wr) arr_me3_f_global_v_E0_i_e_0069 <= out;
   if (mem_addr_wr == 198 && mem_wr) arr_me3_f_global_v_E0_i_e_0070 <= out;
   if (mem_addr_wr == 199 && mem_wr) arr_me3_f_global_v_E0_i_e_0071 <= out;
   if (mem_addr_wr == 200 && mem_wr) arr_me3_f_global_v_E0_i_e_0072 <= out;
   if (mem_addr_wr == 201 && mem_wr) arr_me3_f_global_v_E0_i_e_0073 <= out;
   if (mem_addr_wr == 202 && mem_wr) arr_me3_f_global_v_E0_i_e_0074 <= out;
   if (mem_addr_wr == 203 && mem_wr) arr_me3_f_global_v_E0_i_e_0075 <= out;
   if (mem_addr_wr == 204 && mem_wr) arr_me3_f_global_v_E0_i_e_0076 <= out;
   if (mem_addr_wr == 205 && mem_wr) arr_me3_f_global_v_E0_i_e_0077 <= out;
   if (mem_addr_wr == 206 && mem_wr) arr_me3_f_global_v_E0_i_e_0078 <= out;
   if (mem_addr_wr == 207 && mem_wr) arr_me3_f_global_v_E0_i_e_0079 <= out;
   if (mem_addr_wr == 208 && mem_wr) arr_me3_f_global_v_E0_i_e_0080 <= out;
   if (mem_addr_wr == 209 && mem_wr) arr_me3_f_global_v_E0_i_e_0081 <= out;
   if (mem_addr_wr == 210 && mem_wr) arr_me3_f_global_v_E0_i_e_0082 <= out;
   if (mem_addr_wr == 211 && mem_wr) arr_me3_f_global_v_E0_i_e_0083 <= out;
   if (mem_addr_wr == 212 && mem_wr) arr_me3_f_global_v_E0_i_e_0084 <= out;
   if (mem_addr_wr == 213 && mem_wr) arr_me3_f_global_v_E0_i_e_0085 <= out;
   if (mem_addr_wr == 214 && mem_wr) arr_me3_f_global_v_E0_i_e_0086 <= out;
   if (mem_addr_wr == 215 && mem_wr) arr_me3_f_global_v_E0_i_e_0087 <= out;
   if (mem_addr_wr == 216 && mem_wr) arr_me3_f_global_v_E0_i_e_0088 <= out;
   if (mem_addr_wr == 217 && mem_wr) arr_me3_f_global_v_E0_i_e_0089 <= out;
   if (mem_addr_wr == 218 && mem_wr) arr_me3_f_global_v_E0_i_e_0090 <= out;
   if (mem_addr_wr == 219 && mem_wr) arr_me3_f_global_v_E0_i_e_0091 <= out;
   if (mem_addr_wr == 220 && mem_wr) arr_me3_f_global_v_E0_i_e_0092 <= out;
   if (mem_addr_wr == 221 && mem_wr) arr_me3_f_global_v_E0_i_e_0093 <= out;
   if (mem_addr_wr == 222 && mem_wr) arr_me3_f_global_v_E0_i_e_0094 <= out;
   if (mem_addr_wr == 223 && mem_wr) arr_me3_f_global_v_E0_i_e_0095 <= out;
   if (mem_addr_wr == 224 && mem_wr) arr_me3_f_global_v_E0_i_e_0096 <= out;
   if (mem_addr_wr == 225 && mem_wr) arr_me3_f_global_v_E0_i_e_0097 <= out;
   if (mem_addr_wr == 226 && mem_wr) arr_me3_f_global_v_E0_i_e_0098 <= out;
   if (mem_addr_wr == 227 && mem_wr) arr_me3_f_global_v_E0_i_e_0099 <= out;
   if (mem_addr_wr == 228 && mem_wr) arr_me3_f_global_v_E0_i_e_0100 <= out;
   if (mem_addr_wr == 229 && mem_wr) arr_me3_f_global_v_E0_i_e_0101 <= out;
   if (mem_addr_wr == 230 && mem_wr) arr_me3_f_global_v_E0_i_e_0102 <= out;
   if (mem_addr_wr == 231 && mem_wr) arr_me3_f_global_v_E0_i_e_0103 <= out;
   if (mem_addr_wr == 232 && mem_wr) arr_me3_f_global_v_E0_i_e_0104 <= out;
   if (mem_addr_wr == 233 && mem_wr) arr_me3_f_global_v_E0_i_e_0105 <= out;
   if (mem_addr_wr == 234 && mem_wr) arr_me3_f_global_v_E0_i_e_0106 <= out;
   if (mem_addr_wr == 235 && mem_wr) arr_me3_f_global_v_E0_i_e_0107 <= out;
   if (mem_addr_wr == 236 && mem_wr) arr_me3_f_global_v_E0_i_e_0108 <= out;
   if (mem_addr_wr == 237 && mem_wr) arr_me3_f_global_v_E0_i_e_0109 <= out;
   if (mem_addr_wr == 238 && mem_wr) arr_me3_f_global_v_E0_i_e_0110 <= out;
   if (mem_addr_wr == 239 && mem_wr) arr_me3_f_global_v_E0_i_e_0111 <= out;
   if (mem_addr_wr == 240 && mem_wr) arr_me3_f_global_v_E0_i_e_0112 <= out;
   if (mem_addr_wr == 241 && mem_wr) arr_me3_f_global_v_E0_i_e_0113 <= out;
   if (mem_addr_wr == 242 && mem_wr) arr_me3_f_global_v_E0_i_e_0114 <= out;
   if (mem_addr_wr == 243 && mem_wr) arr_me3_f_global_v_E0_i_e_0115 <= out;
   if (mem_addr_wr == 244 && mem_wr) arr_me3_f_global_v_E0_i_e_0116 <= out;
   if (mem_addr_wr == 245 && mem_wr) arr_me3_f_global_v_E0_i_e_0117 <= out;
   if (mem_addr_wr == 246 && mem_wr) arr_me3_f_global_v_E0_i_e_0118 <= out;
   if (mem_addr_wr == 247 && mem_wr) arr_me3_f_global_v_E0_i_e_0119 <= out;
   if (mem_addr_wr == 248 && mem_wr) arr_me3_f_global_v_E0_i_e_0120 <= out;
   if (mem_addr_wr == 249 && mem_wr) arr_me3_f_global_v_E0_i_e_0121 <= out;
   if (mem_addr_wr == 250 && mem_wr) arr_me3_f_global_v_E0_i_e_0122 <= out;
   if (mem_addr_wr == 251 && mem_wr) arr_me3_f_global_v_E0_i_e_0123 <= out;
   if (mem_addr_wr == 252 && mem_wr) arr_me3_f_global_v_E0_i_e_0124 <= out;
   if (mem_addr_wr == 253 && mem_wr) arr_me3_f_global_v_E0_i_e_0125 <= out;
   if (mem_addr_wr == 254 && mem_wr) arr_me3_f_global_v_E0_i_e_0126 <= out;
   if (mem_addr_wr == 255 && mem_wr) arr_me3_f_global_v_E0_i_e_0127 <= out;
   if (mem_addr_wr == 256 && mem_wr) arr_me3_f_global_v_wpv_e_0000 <= out;
   if (mem_addr_wr == 257 && mem_wr) arr_me3_f_global_v_wpv_e_0001 <= out;
   if (mem_addr_wr == 258 && mem_wr) arr_me3_f_global_v_wpv_e_0002 <= out;
   if (mem_addr_wr == 259 && mem_wr) arr_me3_f_global_v_wpv_e_0003 <= out;
   if (mem_addr_wr == 260 && mem_wr) arr_me3_f_global_v_wpv_e_0004 <= out;
   if (mem_addr_wr == 261 && mem_wr) arr_me3_f_global_v_wpv_e_0005 <= out;
   if (mem_addr_wr == 262 && mem_wr) arr_me3_f_global_v_wpv_e_0006 <= out;
   if (mem_addr_wr == 263 && mem_wr) arr_me3_f_global_v_wpv_e_0007 <= out;
   if (mem_addr_wr == 264 && mem_wr) arr_me3_f_global_v_wpv_e_0008 <= out;
   if (mem_addr_wr == 265 && mem_wr) arr_me3_f_global_v_wpv_e_0009 <= out;
   if (mem_addr_wr == 266 && mem_wr) arr_me3_f_global_v_wpv_e_0010 <= out;
   if (mem_addr_wr == 267 && mem_wr) arr_me3_f_global_v_wpv_e_0011 <= out;
   if (mem_addr_wr == 268 && mem_wr) arr_me3_f_global_v_wpv_e_0012 <= out;
   if (mem_addr_wr == 269 && mem_wr) arr_me3_f_global_v_wpv_e_0013 <= out;
   if (mem_addr_wr == 270 && mem_wr) arr_me3_f_global_v_wpv_e_0014 <= out;
   if (mem_addr_wr == 271 && mem_wr) arr_me3_f_global_v_wpv_e_0015 <= out;
   if (mem_addr_wr == 272 && mem_wr) arr_me3_f_global_v_wpv_e_0016 <= out;
   if (mem_addr_wr == 273 && mem_wr) arr_me3_f_global_v_wpv_e_0017 <= out;
   if (mem_addr_wr == 274 && mem_wr) arr_me3_f_global_v_wpv_e_0018 <= out;
   if (mem_addr_wr == 275 && mem_wr) arr_me3_f_global_v_wpv_e_0019 <= out;
   if (mem_addr_wr == 276 && mem_wr) arr_me3_f_global_v_wpv_e_0020 <= out;
   if (mem_addr_wr == 277 && mem_wr) arr_me3_f_global_v_wpv_e_0021 <= out;
   if (mem_addr_wr == 278 && mem_wr) arr_me3_f_global_v_wpv_e_0022 <= out;
   if (mem_addr_wr == 279 && mem_wr) arr_me3_f_global_v_wpv_e_0023 <= out;
   if (mem_addr_wr == 280 && mem_wr) arr_me3_f_global_v_wpv_e_0024 <= out;
   if (mem_addr_wr == 281 && mem_wr) arr_me3_f_global_v_wpv_e_0025 <= out;
   if (mem_addr_wr == 282 && mem_wr) arr_me3_f_global_v_wpv_e_0026 <= out;
   if (mem_addr_wr == 283 && mem_wr) arr_me3_f_global_v_wpv_e_0027 <= out;
   if (mem_addr_wr == 284 && mem_wr) arr_me3_f_global_v_wpv_e_0028 <= out;
   if (mem_addr_wr == 285 && mem_wr) arr_me3_f_global_v_wpv_e_0029 <= out;
   if (mem_addr_wr == 286 && mem_wr) arr_me3_f_global_v_wpv_e_0030 <= out;
   if (mem_addr_wr == 287 && mem_wr) arr_me3_f_global_v_wpv_e_0031 <= out;
   if (mem_addr_wr == 288 && mem_wr) arr_me3_f_global_v_wpv_e_0032 <= out;
   if (mem_addr_wr == 289 && mem_wr) arr_me3_f_global_v_wpv_e_0033 <= out;
   if (mem_addr_wr == 290 && mem_wr) arr_me3_f_global_v_wpv_e_0034 <= out;
   if (mem_addr_wr == 291 && mem_wr) arr_me3_f_global_v_wpv_e_0035 <= out;
   if (mem_addr_wr == 292 && mem_wr) arr_me3_f_global_v_wpv_e_0036 <= out;
   if (mem_addr_wr == 293 && mem_wr) arr_me3_f_global_v_wpv_e_0037 <= out;
   if (mem_addr_wr == 294 && mem_wr) arr_me3_f_global_v_wpv_e_0038 <= out;
   if (mem_addr_wr == 295 && mem_wr) arr_me3_f_global_v_wpv_e_0039 <= out;
   if (mem_addr_wr == 296 && mem_wr) arr_me3_f_global_v_wpv_e_0040 <= out;
   if (mem_addr_wr == 297 && mem_wr) arr_me3_f_global_v_wpv_e_0041 <= out;
   if (mem_addr_wr == 298 && mem_wr) arr_me3_f_global_v_wpv_e_0042 <= out;
   if (mem_addr_wr == 299 && mem_wr) arr_me3_f_global_v_wpv_e_0043 <= out;
   if (mem_addr_wr == 300 && mem_wr) arr_me3_f_global_v_wpv_e_0044 <= out;
   if (mem_addr_wr == 301 && mem_wr) arr_me3_f_global_v_wpv_e_0045 <= out;
   if (mem_addr_wr == 302 && mem_wr) arr_me3_f_global_v_wpv_e_0046 <= out;
   if (mem_addr_wr == 303 && mem_wr) arr_me3_f_global_v_wpv_e_0047 <= out;
   if (mem_addr_wr == 304 && mem_wr) arr_me3_f_global_v_wpv_e_0048 <= out;
   if (mem_addr_wr == 305 && mem_wr) arr_me3_f_global_v_wpv_e_0049 <= out;
   if (mem_addr_wr == 306 && mem_wr) arr_me3_f_global_v_wpv_e_0050 <= out;
   if (mem_addr_wr == 307 && mem_wr) arr_me3_f_global_v_wpv_e_0051 <= out;
   if (mem_addr_wr == 308 && mem_wr) arr_me3_f_global_v_wpv_e_0052 <= out;
   if (mem_addr_wr == 309 && mem_wr) arr_me3_f_global_v_wpv_e_0053 <= out;
   if (mem_addr_wr == 310 && mem_wr) arr_me3_f_global_v_wpv_e_0054 <= out;
   if (mem_addr_wr == 311 && mem_wr) arr_me3_f_global_v_wpv_e_0055 <= out;
   if (mem_addr_wr == 312 && mem_wr) arr_me3_f_global_v_wpv_e_0056 <= out;
   if (mem_addr_wr == 313 && mem_wr) arr_me3_f_global_v_wpv_e_0057 <= out;
   if (mem_addr_wr == 314 && mem_wr) arr_me3_f_global_v_wpv_e_0058 <= out;
   if (mem_addr_wr == 315 && mem_wr) arr_me3_f_global_v_wpv_e_0059 <= out;
   if (mem_addr_wr == 316 && mem_wr) arr_me3_f_global_v_wpv_e_0060 <= out;
   if (mem_addr_wr == 317 && mem_wr) arr_me3_f_global_v_wpv_e_0061 <= out;
   if (mem_addr_wr == 318 && mem_wr) arr_me3_f_global_v_wpv_e_0062 <= out;
   if (mem_addr_wr == 319 && mem_wr) arr_me3_f_global_v_wpv_e_0063 <= out;
   if (mem_addr_wr == 320 && mem_wr) arr_me3_f_global_v_wpv_i_e_0000 <= out;
   if (mem_addr_wr == 321 && mem_wr) arr_me3_f_global_v_wpv_i_e_0001 <= out;
   if (mem_addr_wr == 322 && mem_wr) arr_me3_f_global_v_wpv_i_e_0002 <= out;
   if (mem_addr_wr == 323 && mem_wr) arr_me3_f_global_v_wpv_i_e_0003 <= out;
   if (mem_addr_wr == 324 && mem_wr) arr_me3_f_global_v_wpv_i_e_0004 <= out;
   if (mem_addr_wr == 325 && mem_wr) arr_me3_f_global_v_wpv_i_e_0005 <= out;
   if (mem_addr_wr == 326 && mem_wr) arr_me3_f_global_v_wpv_i_e_0006 <= out;
   if (mem_addr_wr == 327 && mem_wr) arr_me3_f_global_v_wpv_i_e_0007 <= out;
   if (mem_addr_wr == 328 && mem_wr) arr_me3_f_global_v_wpv_i_e_0008 <= out;
   if (mem_addr_wr == 329 && mem_wr) arr_me3_f_global_v_wpv_i_e_0009 <= out;
   if (mem_addr_wr == 330 && mem_wr) arr_me3_f_global_v_wpv_i_e_0010 <= out;
   if (mem_addr_wr == 331 && mem_wr) arr_me3_f_global_v_wpv_i_e_0011 <= out;
   if (mem_addr_wr == 332 && mem_wr) arr_me3_f_global_v_wpv_i_e_0012 <= out;
   if (mem_addr_wr == 333 && mem_wr) arr_me3_f_global_v_wpv_i_e_0013 <= out;
   if (mem_addr_wr == 334 && mem_wr) arr_me3_f_global_v_wpv_i_e_0014 <= out;
   if (mem_addr_wr == 335 && mem_wr) arr_me3_f_global_v_wpv_i_e_0015 <= out;
   if (mem_addr_wr == 336 && mem_wr) arr_me3_f_global_v_wpv_i_e_0016 <= out;
   if (mem_addr_wr == 337 && mem_wr) arr_me3_f_global_v_wpv_i_e_0017 <= out;
   if (mem_addr_wr == 338 && mem_wr) arr_me3_f_global_v_wpv_i_e_0018 <= out;
   if (mem_addr_wr == 339 && mem_wr) arr_me3_f_global_v_wpv_i_e_0019 <= out;
   if (mem_addr_wr == 340 && mem_wr) arr_me3_f_global_v_wpv_i_e_0020 <= out;
   if (mem_addr_wr == 341 && mem_wr) arr_me3_f_global_v_wpv_i_e_0021 <= out;
   if (mem_addr_wr == 342 && mem_wr) arr_me3_f_global_v_wpv_i_e_0022 <= out;
   if (mem_addr_wr == 343 && mem_wr) arr_me3_f_global_v_wpv_i_e_0023 <= out;
   if (mem_addr_wr == 344 && mem_wr) arr_me3_f_global_v_wpv_i_e_0024 <= out;
   if (mem_addr_wr == 345 && mem_wr) arr_me3_f_global_v_wpv_i_e_0025 <= out;
   if (mem_addr_wr == 346 && mem_wr) arr_me3_f_global_v_wpv_i_e_0026 <= out;
   if (mem_addr_wr == 347 && mem_wr) arr_me3_f_global_v_wpv_i_e_0027 <= out;
   if (mem_addr_wr == 348 && mem_wr) arr_me3_f_global_v_wpv_i_e_0028 <= out;
   if (mem_addr_wr == 349 && mem_wr) arr_me3_f_global_v_wpv_i_e_0029 <= out;
   if (mem_addr_wr == 350 && mem_wr) arr_me3_f_global_v_wpv_i_e_0030 <= out;
   if (mem_addr_wr == 351 && mem_wr) arr_me3_f_global_v_wpv_i_e_0031 <= out;
   if (mem_addr_wr == 352 && mem_wr) arr_me3_f_global_v_wpv_i_e_0032 <= out;
   if (mem_addr_wr == 353 && mem_wr) arr_me3_f_global_v_wpv_i_e_0033 <= out;
   if (mem_addr_wr == 354 && mem_wr) arr_me3_f_global_v_wpv_i_e_0034 <= out;
   if (mem_addr_wr == 355 && mem_wr) arr_me3_f_global_v_wpv_i_e_0035 <= out;
   if (mem_addr_wr == 356 && mem_wr) arr_me3_f_global_v_wpv_i_e_0036 <= out;
   if (mem_addr_wr == 357 && mem_wr) arr_me3_f_global_v_wpv_i_e_0037 <= out;
   if (mem_addr_wr == 358 && mem_wr) arr_me3_f_global_v_wpv_i_e_0038 <= out;
   if (mem_addr_wr == 359 && mem_wr) arr_me3_f_global_v_wpv_i_e_0039 <= out;
   if (mem_addr_wr == 360 && mem_wr) arr_me3_f_global_v_wpv_i_e_0040 <= out;
   if (mem_addr_wr == 361 && mem_wr) arr_me3_f_global_v_wpv_i_e_0041 <= out;
   if (mem_addr_wr == 362 && mem_wr) arr_me3_f_global_v_wpv_i_e_0042 <= out;
   if (mem_addr_wr == 363 && mem_wr) arr_me3_f_global_v_wpv_i_e_0043 <= out;
   if (mem_addr_wr == 364 && mem_wr) arr_me3_f_global_v_wpv_i_e_0044 <= out;
   if (mem_addr_wr == 365 && mem_wr) arr_me3_f_global_v_wpv_i_e_0045 <= out;
   if (mem_addr_wr == 366 && mem_wr) arr_me3_f_global_v_wpv_i_e_0046 <= out;
   if (mem_addr_wr == 367 && mem_wr) arr_me3_f_global_v_wpv_i_e_0047 <= out;
   if (mem_addr_wr == 368 && mem_wr) arr_me3_f_global_v_wpv_i_e_0048 <= out;
   if (mem_addr_wr == 369 && mem_wr) arr_me3_f_global_v_wpv_i_e_0049 <= out;
   if (mem_addr_wr == 370 && mem_wr) arr_me3_f_global_v_wpv_i_e_0050 <= out;
   if (mem_addr_wr == 371 && mem_wr) arr_me3_f_global_v_wpv_i_e_0051 <= out;
   if (mem_addr_wr == 372 && mem_wr) arr_me3_f_global_v_wpv_i_e_0052 <= out;
   if (mem_addr_wr == 373 && mem_wr) arr_me3_f_global_v_wpv_i_e_0053 <= out;
   if (mem_addr_wr == 374 && mem_wr) arr_me3_f_global_v_wpv_i_e_0054 <= out;
   if (mem_addr_wr == 375 && mem_wr) arr_me3_f_global_v_wpv_i_e_0055 <= out;
   if (mem_addr_wr == 376 && mem_wr) arr_me3_f_global_v_wpv_i_e_0056 <= out;
   if (mem_addr_wr == 377 && mem_wr) arr_me3_f_global_v_wpv_i_e_0057 <= out;
   if (mem_addr_wr == 378 && mem_wr) arr_me3_f_global_v_wpv_i_e_0058 <= out;
   if (mem_addr_wr == 379 && mem_wr) arr_me3_f_global_v_wpv_i_e_0059 <= out;
   if (mem_addr_wr == 380 && mem_wr) arr_me3_f_global_v_wpv_i_e_0060 <= out;
   if (mem_addr_wr == 381 && mem_wr) arr_me3_f_global_v_wpv_i_e_0061 <= out;
   if (mem_addr_wr == 382 && mem_wr) arr_me3_f_global_v_wpv_i_e_0062 <= out;
   if (mem_addr_wr == 383 && mem_wr) arr_me3_f_global_v_wpv_i_e_0063 <= out;
   if (mem_addr_wr == 403 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0000 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 404 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0001 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 405 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0002 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 406 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0003 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 407 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0004 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 408 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0005 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 409 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0006 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 410 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0007 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 411 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0008 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 412 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0009 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 413 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0010 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 414 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0011 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 415 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0012 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 416 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0013 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 417 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0014 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 418 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0015 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 419 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0016 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 420 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0017 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 421 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0018 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 422 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0019 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 423 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0020 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 424 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0021 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 425 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0022 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 426 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0023 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 427 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0024 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 428 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0025 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 429 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0026 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 430 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0027 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 431 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0028 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 432 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0029 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 433 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0030 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 434 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0031 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 435 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0032 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 436 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0033 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 437 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0034 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 438 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0035 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 439 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0036 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 440 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0037 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 441 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0038 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 442 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0039 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 443 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0040 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 444 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0041 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 445 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0042 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 446 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0043 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 447 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0044 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 448 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0045 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 449 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0046 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 450 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0047 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 451 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0048 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 452 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0049 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 453 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0050 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 454 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0051 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 455 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0052 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 456 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0053 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 457 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0054 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 458 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0055 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 459 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0056 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 460 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0057 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 461 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0058 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 462 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0059 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 463 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0060 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 464 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0061 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 465 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0062 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 466 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0063 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 467 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0064 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 468 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0065 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 469 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0066 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 470 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0067 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 471 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0068 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 472 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0069 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 473 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0070 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 474 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0071 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 475 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0072 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 476 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0073 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 477 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0074 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 478 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0075 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 479 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0076 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 480 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0077 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 481 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0078 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 482 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0079 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 483 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0080 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 484 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0081 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 485 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0082 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 486 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0083 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 487 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0084 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 488 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0085 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 489 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0086 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 490 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0087 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 491 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0088 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 492 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0089 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 493 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0090 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 494 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0091 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 495 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0092 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 496 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0093 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 497 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0094 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 498 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0095 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 499 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0096 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 500 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0097 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 501 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0098 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 502 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0099 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 503 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0100 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 504 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0101 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 505 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0102 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 506 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0103 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 507 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0104 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 508 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0105 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 509 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0106 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 510 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0107 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 511 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0108 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 512 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0109 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 513 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0110 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 514 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0111 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 515 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0112 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 516 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0113 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 517 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0114 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 518 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0115 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 519 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0116 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 520 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0117 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 521 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0118 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 522 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0119 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 523 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0120 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 524 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0121 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 525 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0122 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 526 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0123 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 527 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0124 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 528 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0125 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 529 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0126 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 530 && mem_wr) arr_me2_f_main_v_output_buffer_real_e_0127 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 531 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0000 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 532 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0001 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 533 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0002 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 534 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0003 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 535 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0004 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 536 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0005 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 537 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0006 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 538 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0007 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 539 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0008 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 540 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0009 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 541 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0010 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 542 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0011 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 543 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0012 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 544 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0013 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 545 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0014 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 546 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0015 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 547 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0016 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 548 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0017 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 549 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0018 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 550 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0019 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 551 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0020 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 552 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0021 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 553 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0022 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 554 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0023 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 555 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0024 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 556 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0025 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 557 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0026 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 558 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0027 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 559 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0028 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 560 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0029 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 561 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0030 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 562 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0031 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 563 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0032 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 564 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0033 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 565 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0034 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 566 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0035 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 567 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0036 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 568 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0037 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 569 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0038 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 570 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0039 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 571 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0040 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 572 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0041 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 573 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0042 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 574 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0043 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 575 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0044 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 576 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0045 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 577 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0046 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 578 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0047 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 579 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0048 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 580 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0049 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 581 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0050 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 582 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0051 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 583 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0052 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 584 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0053 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 585 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0054 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 586 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0055 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 587 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0056 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 588 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0057 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 589 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0058 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 590 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0059 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 591 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0060 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 592 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0061 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 593 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0062 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 594 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0063 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 595 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0064 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 596 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0065 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 597 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0066 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 598 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0067 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 599 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0068 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 600 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0069 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 601 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0070 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 602 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0071 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 603 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0072 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 604 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0073 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 605 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0074 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 606 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0075 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 607 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0076 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 608 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0077 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 609 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0078 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 610 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0079 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 611 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0080 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 612 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0081 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 613 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0082 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 614 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0083 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 615 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0084 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 616 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0085 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 617 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0086 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 618 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0087 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 619 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0088 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 620 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0089 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 621 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0090 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 622 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0091 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 623 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0092 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 624 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0093 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 625 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0094 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 626 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0095 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 627 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0096 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 628 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0097 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 629 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0098 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 630 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0099 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 631 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0100 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 632 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0101 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 633 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0102 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 634 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0103 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 635 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0104 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 636 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0105 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 637 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0106 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 638 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0107 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 639 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0108 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 640 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0109 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 641 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0110 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 642 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0111 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 643 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0112 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 644 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0113 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 645 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0114 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 646 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0115 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 647 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0116 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 648 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0117 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 649 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0118 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 650 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0119 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 651 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0120 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 652 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0121 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 653 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0122 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 654 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0123 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 655 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0124 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 656 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0125 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 657 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0126 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 658 && mem_wr) arr_me2_f_main_v_output_buffer_imag_e_0127 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 659 && mem_wr) arr_me2_f_main_v_buffer_e_0000 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 660 && mem_wr) arr_me2_f_main_v_buffer_e_0001 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 661 && mem_wr) arr_me2_f_main_v_buffer_e_0002 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 662 && mem_wr) arr_me2_f_main_v_buffer_e_0003 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 663 && mem_wr) arr_me2_f_main_v_buffer_e_0004 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 664 && mem_wr) arr_me2_f_main_v_buffer_e_0005 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 665 && mem_wr) arr_me2_f_main_v_buffer_e_0006 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 666 && mem_wr) arr_me2_f_main_v_buffer_e_0007 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 667 && mem_wr) arr_me2_f_main_v_buffer_e_0008 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 668 && mem_wr) arr_me2_f_main_v_buffer_e_0009 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 669 && mem_wr) arr_me2_f_main_v_buffer_e_0010 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 670 && mem_wr) arr_me2_f_main_v_buffer_e_0011 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 671 && mem_wr) arr_me2_f_main_v_buffer_e_0012 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 672 && mem_wr) arr_me2_f_main_v_buffer_e_0013 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 673 && mem_wr) arr_me2_f_main_v_buffer_e_0014 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 674 && mem_wr) arr_me2_f_main_v_buffer_e_0015 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 675 && mem_wr) arr_me2_f_main_v_buffer_e_0016 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 676 && mem_wr) arr_me2_f_main_v_buffer_e_0017 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 677 && mem_wr) arr_me2_f_main_v_buffer_e_0018 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 678 && mem_wr) arr_me2_f_main_v_buffer_e_0019 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 679 && mem_wr) arr_me2_f_main_v_buffer_e_0020 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 680 && mem_wr) arr_me2_f_main_v_buffer_e_0021 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 681 && mem_wr) arr_me2_f_main_v_buffer_e_0022 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 682 && mem_wr) arr_me2_f_main_v_buffer_e_0023 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 683 && mem_wr) arr_me2_f_main_v_buffer_e_0024 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 684 && mem_wr) arr_me2_f_main_v_buffer_e_0025 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 685 && mem_wr) arr_me2_f_main_v_buffer_e_0026 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 686 && mem_wr) arr_me2_f_main_v_buffer_e_0027 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 687 && mem_wr) arr_me2_f_main_v_buffer_e_0028 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 688 && mem_wr) arr_me2_f_main_v_buffer_e_0029 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 689 && mem_wr) arr_me2_f_main_v_buffer_e_0030 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 690 && mem_wr) arr_me2_f_main_v_buffer_e_0031 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 691 && mem_wr) arr_me2_f_main_v_buffer_e_0032 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 692 && mem_wr) arr_me2_f_main_v_buffer_e_0033 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 693 && mem_wr) arr_me2_f_main_v_buffer_e_0034 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 694 && mem_wr) arr_me2_f_main_v_buffer_e_0035 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 695 && mem_wr) arr_me2_f_main_v_buffer_e_0036 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 696 && mem_wr) arr_me2_f_main_v_buffer_e_0037 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 697 && mem_wr) arr_me2_f_main_v_buffer_e_0038 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 698 && mem_wr) arr_me2_f_main_v_buffer_e_0039 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 699 && mem_wr) arr_me2_f_main_v_buffer_e_0040 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 700 && mem_wr) arr_me2_f_main_v_buffer_e_0041 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 701 && mem_wr) arr_me2_f_main_v_buffer_e_0042 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 702 && mem_wr) arr_me2_f_main_v_buffer_e_0043 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 703 && mem_wr) arr_me2_f_main_v_buffer_e_0044 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 704 && mem_wr) arr_me2_f_main_v_buffer_e_0045 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 705 && mem_wr) arr_me2_f_main_v_buffer_e_0046 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 706 && mem_wr) arr_me2_f_main_v_buffer_e_0047 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 707 && mem_wr) arr_me2_f_main_v_buffer_e_0048 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 708 && mem_wr) arr_me2_f_main_v_buffer_e_0049 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 709 && mem_wr) arr_me2_f_main_v_buffer_e_0050 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 710 && mem_wr) arr_me2_f_main_v_buffer_e_0051 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 711 && mem_wr) arr_me2_f_main_v_buffer_e_0052 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 712 && mem_wr) arr_me2_f_main_v_buffer_e_0053 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 713 && mem_wr) arr_me2_f_main_v_buffer_e_0054 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 714 && mem_wr) arr_me2_f_main_v_buffer_e_0055 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 715 && mem_wr) arr_me2_f_main_v_buffer_e_0056 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 716 && mem_wr) arr_me2_f_main_v_buffer_e_0057 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 717 && mem_wr) arr_me2_f_main_v_buffer_e_0058 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 718 && mem_wr) arr_me2_f_main_v_buffer_e_0059 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 719 && mem_wr) arr_me2_f_main_v_buffer_e_0060 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 720 && mem_wr) arr_me2_f_main_v_buffer_e_0061 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 721 && mem_wr) arr_me2_f_main_v_buffer_e_0062 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 722 && mem_wr) arr_me2_f_main_v_buffer_e_0063 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 723 && mem_wr) arr_me2_f_main_v_buffer_e_0064 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 724 && mem_wr) arr_me2_f_main_v_buffer_e_0065 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 725 && mem_wr) arr_me2_f_main_v_buffer_e_0066 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 726 && mem_wr) arr_me2_f_main_v_buffer_e_0067 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 727 && mem_wr) arr_me2_f_main_v_buffer_e_0068 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 728 && mem_wr) arr_me2_f_main_v_buffer_e_0069 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 729 && mem_wr) arr_me2_f_main_v_buffer_e_0070 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 730 && mem_wr) arr_me2_f_main_v_buffer_e_0071 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 731 && mem_wr) arr_me2_f_main_v_buffer_e_0072 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 732 && mem_wr) arr_me2_f_main_v_buffer_e_0073 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 733 && mem_wr) arr_me2_f_main_v_buffer_e_0074 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 734 && mem_wr) arr_me2_f_main_v_buffer_e_0075 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 735 && mem_wr) arr_me2_f_main_v_buffer_e_0076 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 736 && mem_wr) arr_me2_f_main_v_buffer_e_0077 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 737 && mem_wr) arr_me2_f_main_v_buffer_e_0078 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 738 && mem_wr) arr_me2_f_main_v_buffer_e_0079 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 739 && mem_wr) arr_me2_f_main_v_buffer_e_0080 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 740 && mem_wr) arr_me2_f_main_v_buffer_e_0081 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 741 && mem_wr) arr_me2_f_main_v_buffer_e_0082 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 742 && mem_wr) arr_me2_f_main_v_buffer_e_0083 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 743 && mem_wr) arr_me2_f_main_v_buffer_e_0084 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 744 && mem_wr) arr_me2_f_main_v_buffer_e_0085 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 745 && mem_wr) arr_me2_f_main_v_buffer_e_0086 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 746 && mem_wr) arr_me2_f_main_v_buffer_e_0087 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 747 && mem_wr) arr_me2_f_main_v_buffer_e_0088 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 748 && mem_wr) arr_me2_f_main_v_buffer_e_0089 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 749 && mem_wr) arr_me2_f_main_v_buffer_e_0090 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 750 && mem_wr) arr_me2_f_main_v_buffer_e_0091 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 751 && mem_wr) arr_me2_f_main_v_buffer_e_0092 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 752 && mem_wr) arr_me2_f_main_v_buffer_e_0093 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 753 && mem_wr) arr_me2_f_main_v_buffer_e_0094 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 754 && mem_wr) arr_me2_f_main_v_buffer_e_0095 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 755 && mem_wr) arr_me2_f_main_v_buffer_e_0096 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 756 && mem_wr) arr_me2_f_main_v_buffer_e_0097 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 757 && mem_wr) arr_me2_f_main_v_buffer_e_0098 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 758 && mem_wr) arr_me2_f_main_v_buffer_e_0099 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 759 && mem_wr) arr_me2_f_main_v_buffer_e_0100 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 760 && mem_wr) arr_me2_f_main_v_buffer_e_0101 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 761 && mem_wr) arr_me2_f_main_v_buffer_e_0102 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 762 && mem_wr) arr_me2_f_main_v_buffer_e_0103 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 763 && mem_wr) arr_me2_f_main_v_buffer_e_0104 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 764 && mem_wr) arr_me2_f_main_v_buffer_e_0105 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 765 && mem_wr) arr_me2_f_main_v_buffer_e_0106 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 766 && mem_wr) arr_me2_f_main_v_buffer_e_0107 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 767 && mem_wr) arr_me2_f_main_v_buffer_e_0108 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 768 && mem_wr) arr_me2_f_main_v_buffer_e_0109 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 769 && mem_wr) arr_me2_f_main_v_buffer_e_0110 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 770 && mem_wr) arr_me2_f_main_v_buffer_e_0111 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 771 && mem_wr) arr_me2_f_main_v_buffer_e_0112 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 772 && mem_wr) arr_me2_f_main_v_buffer_e_0113 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 773 && mem_wr) arr_me2_f_main_v_buffer_e_0114 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 774 && mem_wr) arr_me2_f_main_v_buffer_e_0115 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 775 && mem_wr) arr_me2_f_main_v_buffer_e_0116 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 776 && mem_wr) arr_me2_f_main_v_buffer_e_0117 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 777 && mem_wr) arr_me2_f_main_v_buffer_e_0118 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 778 && mem_wr) arr_me2_f_main_v_buffer_e_0119 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 779 && mem_wr) arr_me2_f_main_v_buffer_e_0120 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 780 && mem_wr) arr_me2_f_main_v_buffer_e_0121 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 781 && mem_wr) arr_me2_f_main_v_buffer_e_0122 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 782 && mem_wr) arr_me2_f_main_v_buffer_e_0123 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 783 && mem_wr) arr_me2_f_main_v_buffer_e_0124 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 784 && mem_wr) arr_me2_f_main_v_buffer_e_0125 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 785 && mem_wr) arr_me2_f_main_v_buffer_e_0126 <= sm_me2*$pow(2.0,e_me2);
   if (mem_addr_wr == 786 && mem_wr) arr_me2_f_main_v_buffer_e_0127 <= sm_me2*$pow(2.0,e_me2);
end

wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0000 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0000, arr_me3_f_global_v_E0_i_e_0000};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0001 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0001, arr_me3_f_global_v_E0_i_e_0001};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0002 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0002, arr_me3_f_global_v_E0_i_e_0002};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0003 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0003, arr_me3_f_global_v_E0_i_e_0003};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0004 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0004, arr_me3_f_global_v_E0_i_e_0004};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0005 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0005, arr_me3_f_global_v_E0_i_e_0005};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0006 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0006, arr_me3_f_global_v_E0_i_e_0006};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0007 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0007, arr_me3_f_global_v_E0_i_e_0007};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0008 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0008, arr_me3_f_global_v_E0_i_e_0008};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0009 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0009, arr_me3_f_global_v_E0_i_e_0009};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0010 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0010, arr_me3_f_global_v_E0_i_e_0010};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0011 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0011, arr_me3_f_global_v_E0_i_e_0011};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0012 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0012, arr_me3_f_global_v_E0_i_e_0012};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0013 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0013, arr_me3_f_global_v_E0_i_e_0013};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0014 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0014, arr_me3_f_global_v_E0_i_e_0014};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0015 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0015, arr_me3_f_global_v_E0_i_e_0015};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0016 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0016, arr_me3_f_global_v_E0_i_e_0016};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0017 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0017, arr_me3_f_global_v_E0_i_e_0017};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0018 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0018, arr_me3_f_global_v_E0_i_e_0018};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0019 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0019, arr_me3_f_global_v_E0_i_e_0019};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0020 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0020, arr_me3_f_global_v_E0_i_e_0020};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0021 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0021, arr_me3_f_global_v_E0_i_e_0021};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0022 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0022, arr_me3_f_global_v_E0_i_e_0022};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0023 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0023, arr_me3_f_global_v_E0_i_e_0023};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0024 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0024, arr_me3_f_global_v_E0_i_e_0024};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0025 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0025, arr_me3_f_global_v_E0_i_e_0025};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0026 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0026, arr_me3_f_global_v_E0_i_e_0026};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0027 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0027, arr_me3_f_global_v_E0_i_e_0027};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0028 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0028, arr_me3_f_global_v_E0_i_e_0028};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0029 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0029, arr_me3_f_global_v_E0_i_e_0029};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0030 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0030, arr_me3_f_global_v_E0_i_e_0030};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0031 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0031, arr_me3_f_global_v_E0_i_e_0031};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0032 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0032, arr_me3_f_global_v_E0_i_e_0032};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0033 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0033, arr_me3_f_global_v_E0_i_e_0033};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0034 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0034, arr_me3_f_global_v_E0_i_e_0034};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0035 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0035, arr_me3_f_global_v_E0_i_e_0035};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0036 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0036, arr_me3_f_global_v_E0_i_e_0036};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0037 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0037, arr_me3_f_global_v_E0_i_e_0037};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0038 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0038, arr_me3_f_global_v_E0_i_e_0038};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0039 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0039, arr_me3_f_global_v_E0_i_e_0039};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0040 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0040, arr_me3_f_global_v_E0_i_e_0040};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0041 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0041, arr_me3_f_global_v_E0_i_e_0041};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0042 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0042, arr_me3_f_global_v_E0_i_e_0042};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0043 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0043, arr_me3_f_global_v_E0_i_e_0043};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0044 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0044, arr_me3_f_global_v_E0_i_e_0044};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0045 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0045, arr_me3_f_global_v_E0_i_e_0045};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0046 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0046, arr_me3_f_global_v_E0_i_e_0046};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0047 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0047, arr_me3_f_global_v_E0_i_e_0047};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0048 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0048, arr_me3_f_global_v_E0_i_e_0048};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0049 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0049, arr_me3_f_global_v_E0_i_e_0049};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0050 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0050, arr_me3_f_global_v_E0_i_e_0050};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0051 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0051, arr_me3_f_global_v_E0_i_e_0051};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0052 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0052, arr_me3_f_global_v_E0_i_e_0052};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0053 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0053, arr_me3_f_global_v_E0_i_e_0053};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0054 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0054, arr_me3_f_global_v_E0_i_e_0054};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0055 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0055, arr_me3_f_global_v_E0_i_e_0055};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0056 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0056, arr_me3_f_global_v_E0_i_e_0056};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0057 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0057, arr_me3_f_global_v_E0_i_e_0057};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0058 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0058, arr_me3_f_global_v_E0_i_e_0058};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0059 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0059, arr_me3_f_global_v_E0_i_e_0059};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0060 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0060, arr_me3_f_global_v_E0_i_e_0060};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0061 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0061, arr_me3_f_global_v_E0_i_e_0061};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0062 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0062, arr_me3_f_global_v_E0_i_e_0062};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0063 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0063, arr_me3_f_global_v_E0_i_e_0063};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0064 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0064, arr_me3_f_global_v_E0_i_e_0064};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0065 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0065, arr_me3_f_global_v_E0_i_e_0065};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0066 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0066, arr_me3_f_global_v_E0_i_e_0066};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0067 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0067, arr_me3_f_global_v_E0_i_e_0067};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0068 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0068, arr_me3_f_global_v_E0_i_e_0068};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0069 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0069, arr_me3_f_global_v_E0_i_e_0069};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0070 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0070, arr_me3_f_global_v_E0_i_e_0070};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0071 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0071, arr_me3_f_global_v_E0_i_e_0071};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0072 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0072, arr_me3_f_global_v_E0_i_e_0072};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0073 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0073, arr_me3_f_global_v_E0_i_e_0073};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0074 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0074, arr_me3_f_global_v_E0_i_e_0074};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0075 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0075, arr_me3_f_global_v_E0_i_e_0075};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0076 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0076, arr_me3_f_global_v_E0_i_e_0076};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0077 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0077, arr_me3_f_global_v_E0_i_e_0077};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0078 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0078, arr_me3_f_global_v_E0_i_e_0078};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0079 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0079, arr_me3_f_global_v_E0_i_e_0079};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0080 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0080, arr_me3_f_global_v_E0_i_e_0080};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0081 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0081, arr_me3_f_global_v_E0_i_e_0081};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0082 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0082, arr_me3_f_global_v_E0_i_e_0082};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0083 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0083, arr_me3_f_global_v_E0_i_e_0083};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0084 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0084, arr_me3_f_global_v_E0_i_e_0084};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0085 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0085, arr_me3_f_global_v_E0_i_e_0085};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0086 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0086, arr_me3_f_global_v_E0_i_e_0086};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0087 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0087, arr_me3_f_global_v_E0_i_e_0087};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0088 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0088, arr_me3_f_global_v_E0_i_e_0088};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0089 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0089, arr_me3_f_global_v_E0_i_e_0089};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0090 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0090, arr_me3_f_global_v_E0_i_e_0090};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0091 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0091, arr_me3_f_global_v_E0_i_e_0091};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0092 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0092, arr_me3_f_global_v_E0_i_e_0092};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0093 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0093, arr_me3_f_global_v_E0_i_e_0093};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0094 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0094, arr_me3_f_global_v_E0_i_e_0094};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0095 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0095, arr_me3_f_global_v_E0_i_e_0095};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0096 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0096, arr_me3_f_global_v_E0_i_e_0096};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0097 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0097, arr_me3_f_global_v_E0_i_e_0097};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0098 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0098, arr_me3_f_global_v_E0_i_e_0098};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0099 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0099, arr_me3_f_global_v_E0_i_e_0099};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0100 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0100, arr_me3_f_global_v_E0_i_e_0100};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0101 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0101, arr_me3_f_global_v_E0_i_e_0101};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0102 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0102, arr_me3_f_global_v_E0_i_e_0102};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0103 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0103, arr_me3_f_global_v_E0_i_e_0103};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0104 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0104, arr_me3_f_global_v_E0_i_e_0104};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0105 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0105, arr_me3_f_global_v_E0_i_e_0105};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0106 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0106, arr_me3_f_global_v_E0_i_e_0106};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0107 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0107, arr_me3_f_global_v_E0_i_e_0107};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0108 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0108, arr_me3_f_global_v_E0_i_e_0108};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0109 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0109, arr_me3_f_global_v_E0_i_e_0109};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0110 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0110, arr_me3_f_global_v_E0_i_e_0110};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0111 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0111, arr_me3_f_global_v_E0_i_e_0111};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0112 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0112, arr_me3_f_global_v_E0_i_e_0112};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0113 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0113, arr_me3_f_global_v_E0_i_e_0113};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0114 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0114, arr_me3_f_global_v_E0_i_e_0114};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0115 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0115, arr_me3_f_global_v_E0_i_e_0115};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0116 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0116, arr_me3_f_global_v_E0_i_e_0116};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0117 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0117, arr_me3_f_global_v_E0_i_e_0117};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0118 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0118, arr_me3_f_global_v_E0_i_e_0118};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0119 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0119, arr_me3_f_global_v_E0_i_e_0119};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0120 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0120, arr_me3_f_global_v_E0_i_e_0120};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0121 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0121, arr_me3_f_global_v_E0_i_e_0121};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0122 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0122, arr_me3_f_global_v_E0_i_e_0122};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0123 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0123, arr_me3_f_global_v_E0_i_e_0123};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0124 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0124, arr_me3_f_global_v_E0_i_e_0124};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0125 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0125, arr_me3_f_global_v_E0_i_e_0125};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0126 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0126, arr_me3_f_global_v_E0_i_e_0126};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_E0_e_0127 = {8'd23, 8'd8, arr_me3_f_global_v_E0_e_0127, arr_me3_f_global_v_E0_i_e_0127};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_wpv_e_0000 = {8'd23, 8'd8, arr_me3_f_global_v_wpv_e_0000, arr_me3_f_global_v_wpv_i_e_0000};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_wpv_e_0001 = {8'd23, 8'd8, arr_me3_f_global_v_wpv_e_0001, arr_me3_f_global_v_wpv_i_e_0001};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_wpv_e_0002 = {8'd23, 8'd8, arr_me3_f_global_v_wpv_e_0002, arr_me3_f_global_v_wpv_i_e_0002};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_wpv_e_0003 = {8'd23, 8'd8, arr_me3_f_global_v_wpv_e_0003, arr_me3_f_global_v_wpv_i_e_0003};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_wpv_e_0004 = {8'd23, 8'd8, arr_me3_f_global_v_wpv_e_0004, arr_me3_f_global_v_wpv_i_e_0004};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_wpv_e_0005 = {8'd23, 8'd8, arr_me3_f_global_v_wpv_e_0005, arr_me3_f_global_v_wpv_i_e_0005};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_wpv_e_0006 = {8'd23, 8'd8, arr_me3_f_global_v_wpv_e_0006, arr_me3_f_global_v_wpv_i_e_0006};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_wpv_e_0007 = {8'd23, 8'd8, arr_me3_f_global_v_wpv_e_0007, arr_me3_f_global_v_wpv_i_e_0007};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_wpv_e_0008 = {8'd23, 8'd8, arr_me3_f_global_v_wpv_e_0008, arr_me3_f_global_v_wpv_i_e_0008};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_wpv_e_0009 = {8'd23, 8'd8, arr_me3_f_global_v_wpv_e_0009, arr_me3_f_global_v_wpv_i_e_0009};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_wpv_e_0010 = {8'd23, 8'd8, arr_me3_f_global_v_wpv_e_0010, arr_me3_f_global_v_wpv_i_e_0010};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_wpv_e_0011 = {8'd23, 8'd8, arr_me3_f_global_v_wpv_e_0011, arr_me3_f_global_v_wpv_i_e_0011};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_wpv_e_0012 = {8'd23, 8'd8, arr_me3_f_global_v_wpv_e_0012, arr_me3_f_global_v_wpv_i_e_0012};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_wpv_e_0013 = {8'd23, 8'd8, arr_me3_f_global_v_wpv_e_0013, arr_me3_f_global_v_wpv_i_e_0013};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_wpv_e_0014 = {8'd23, 8'd8, arr_me3_f_global_v_wpv_e_0014, arr_me3_f_global_v_wpv_i_e_0014};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_wpv_e_0015 = {8'd23, 8'd8, arr_me3_f_global_v_wpv_e_0015, arr_me3_f_global_v_wpv_i_e_0015};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_wpv_e_0016 = {8'd23, 8'd8, arr_me3_f_global_v_wpv_e_0016, arr_me3_f_global_v_wpv_i_e_0016};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_wpv_e_0017 = {8'd23, 8'd8, arr_me3_f_global_v_wpv_e_0017, arr_me3_f_global_v_wpv_i_e_0017};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_wpv_e_0018 = {8'd23, 8'd8, arr_me3_f_global_v_wpv_e_0018, arr_me3_f_global_v_wpv_i_e_0018};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_wpv_e_0019 = {8'd23, 8'd8, arr_me3_f_global_v_wpv_e_0019, arr_me3_f_global_v_wpv_i_e_0019};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_wpv_e_0020 = {8'd23, 8'd8, arr_me3_f_global_v_wpv_e_0020, arr_me3_f_global_v_wpv_i_e_0020};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_wpv_e_0021 = {8'd23, 8'd8, arr_me3_f_global_v_wpv_e_0021, arr_me3_f_global_v_wpv_i_e_0021};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_wpv_e_0022 = {8'd23, 8'd8, arr_me3_f_global_v_wpv_e_0022, arr_me3_f_global_v_wpv_i_e_0022};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_wpv_e_0023 = {8'd23, 8'd8, arr_me3_f_global_v_wpv_e_0023, arr_me3_f_global_v_wpv_i_e_0023};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_wpv_e_0024 = {8'd23, 8'd8, arr_me3_f_global_v_wpv_e_0024, arr_me3_f_global_v_wpv_i_e_0024};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_wpv_e_0025 = {8'd23, 8'd8, arr_me3_f_global_v_wpv_e_0025, arr_me3_f_global_v_wpv_i_e_0025};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_wpv_e_0026 = {8'd23, 8'd8, arr_me3_f_global_v_wpv_e_0026, arr_me3_f_global_v_wpv_i_e_0026};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_wpv_e_0027 = {8'd23, 8'd8, arr_me3_f_global_v_wpv_e_0027, arr_me3_f_global_v_wpv_i_e_0027};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_wpv_e_0028 = {8'd23, 8'd8, arr_me3_f_global_v_wpv_e_0028, arr_me3_f_global_v_wpv_i_e_0028};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_wpv_e_0029 = {8'd23, 8'd8, arr_me3_f_global_v_wpv_e_0029, arr_me3_f_global_v_wpv_i_e_0029};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_wpv_e_0030 = {8'd23, 8'd8, arr_me3_f_global_v_wpv_e_0030, arr_me3_f_global_v_wpv_i_e_0030};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_wpv_e_0031 = {8'd23, 8'd8, arr_me3_f_global_v_wpv_e_0031, arr_me3_f_global_v_wpv_i_e_0031};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_wpv_e_0032 = {8'd23, 8'd8, arr_me3_f_global_v_wpv_e_0032, arr_me3_f_global_v_wpv_i_e_0032};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_wpv_e_0033 = {8'd23, 8'd8, arr_me3_f_global_v_wpv_e_0033, arr_me3_f_global_v_wpv_i_e_0033};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_wpv_e_0034 = {8'd23, 8'd8, arr_me3_f_global_v_wpv_e_0034, arr_me3_f_global_v_wpv_i_e_0034};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_wpv_e_0035 = {8'd23, 8'd8, arr_me3_f_global_v_wpv_e_0035, arr_me3_f_global_v_wpv_i_e_0035};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_wpv_e_0036 = {8'd23, 8'd8, arr_me3_f_global_v_wpv_e_0036, arr_me3_f_global_v_wpv_i_e_0036};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_wpv_e_0037 = {8'd23, 8'd8, arr_me3_f_global_v_wpv_e_0037, arr_me3_f_global_v_wpv_i_e_0037};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_wpv_e_0038 = {8'd23, 8'd8, arr_me3_f_global_v_wpv_e_0038, arr_me3_f_global_v_wpv_i_e_0038};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_wpv_e_0039 = {8'd23, 8'd8, arr_me3_f_global_v_wpv_e_0039, arr_me3_f_global_v_wpv_i_e_0039};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_wpv_e_0040 = {8'd23, 8'd8, arr_me3_f_global_v_wpv_e_0040, arr_me3_f_global_v_wpv_i_e_0040};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_wpv_e_0041 = {8'd23, 8'd8, arr_me3_f_global_v_wpv_e_0041, arr_me3_f_global_v_wpv_i_e_0041};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_wpv_e_0042 = {8'd23, 8'd8, arr_me3_f_global_v_wpv_e_0042, arr_me3_f_global_v_wpv_i_e_0042};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_wpv_e_0043 = {8'd23, 8'd8, arr_me3_f_global_v_wpv_e_0043, arr_me3_f_global_v_wpv_i_e_0043};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_wpv_e_0044 = {8'd23, 8'd8, arr_me3_f_global_v_wpv_e_0044, arr_me3_f_global_v_wpv_i_e_0044};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_wpv_e_0045 = {8'd23, 8'd8, arr_me3_f_global_v_wpv_e_0045, arr_me3_f_global_v_wpv_i_e_0045};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_wpv_e_0046 = {8'd23, 8'd8, arr_me3_f_global_v_wpv_e_0046, arr_me3_f_global_v_wpv_i_e_0046};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_wpv_e_0047 = {8'd23, 8'd8, arr_me3_f_global_v_wpv_e_0047, arr_me3_f_global_v_wpv_i_e_0047};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_wpv_e_0048 = {8'd23, 8'd8, arr_me3_f_global_v_wpv_e_0048, arr_me3_f_global_v_wpv_i_e_0048};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_wpv_e_0049 = {8'd23, 8'd8, arr_me3_f_global_v_wpv_e_0049, arr_me3_f_global_v_wpv_i_e_0049};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_wpv_e_0050 = {8'd23, 8'd8, arr_me3_f_global_v_wpv_e_0050, arr_me3_f_global_v_wpv_i_e_0050};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_wpv_e_0051 = {8'd23, 8'd8, arr_me3_f_global_v_wpv_e_0051, arr_me3_f_global_v_wpv_i_e_0051};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_wpv_e_0052 = {8'd23, 8'd8, arr_me3_f_global_v_wpv_e_0052, arr_me3_f_global_v_wpv_i_e_0052};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_wpv_e_0053 = {8'd23, 8'd8, arr_me3_f_global_v_wpv_e_0053, arr_me3_f_global_v_wpv_i_e_0053};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_wpv_e_0054 = {8'd23, 8'd8, arr_me3_f_global_v_wpv_e_0054, arr_me3_f_global_v_wpv_i_e_0054};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_wpv_e_0055 = {8'd23, 8'd8, arr_me3_f_global_v_wpv_e_0055, arr_me3_f_global_v_wpv_i_e_0055};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_wpv_e_0056 = {8'd23, 8'd8, arr_me3_f_global_v_wpv_e_0056, arr_me3_f_global_v_wpv_i_e_0056};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_wpv_e_0057 = {8'd23, 8'd8, arr_me3_f_global_v_wpv_e_0057, arr_me3_f_global_v_wpv_i_e_0057};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_wpv_e_0058 = {8'd23, 8'd8, arr_me3_f_global_v_wpv_e_0058, arr_me3_f_global_v_wpv_i_e_0058};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_wpv_e_0059 = {8'd23, 8'd8, arr_me3_f_global_v_wpv_e_0059, arr_me3_f_global_v_wpv_i_e_0059};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_wpv_e_0060 = {8'd23, 8'd8, arr_me3_f_global_v_wpv_e_0060, arr_me3_f_global_v_wpv_i_e_0060};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_wpv_e_0061 = {8'd23, 8'd8, arr_me3_f_global_v_wpv_e_0061, arr_me3_f_global_v_wpv_i_e_0061};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_wpv_e_0062 = {8'd23, 8'd8, arr_me3_f_global_v_wpv_e_0062, arr_me3_f_global_v_wpv_i_e_0062};
wire [16+32*2-1:0] comp_arr_me3_f_global_v_wpv_e_0063 = {8'd23, 8'd8, arr_me3_f_global_v_wpv_e_0063, arr_me3_f_global_v_wpv_i_e_0063};

// instrucoes -----------------------------------------------------------------

reg [31:0] valr1=0;
reg [31:0] valr2=0;
reg [31:0] valr3=0;
reg [31:0] valr4=0;
reg [31:0] valr5=0;
reg [31:0] valr6=0;
reg [31:0] valr7=0;
reg [31:0] valr8=0;
reg [31:0] valr9=0;
reg [31:0] valr10=0;

reg [19:0] min [0:324-1];

reg signed [19:0] linetab =-1;
reg signed [19:0] linetabs=-1;

initial	$readmemb("pc_procTest_00_mem.txt",min);

always @ (posedge clk) begin
if (pc_sim_val < 324) linetab <= min[pc_sim_val];
linetabs <= linetab;   
valr1    <= pc_sim_val;
valr2    <= valr1;
valr3    <= valr2;
valr4    <= valr3;
valr5    <= valr4;
valr6    <= valr5;
valr7    <= valr6;
valr8    <= valr7;
valr9    <= valr8;
valr10   <= valr9;
end

always @ (posedge clk) if (valr10 == 2) begin
   $display("Info: end of program!");
   $finish;
end

`endif

endmodule