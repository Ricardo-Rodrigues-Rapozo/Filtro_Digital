`timescale 1ns/1ps

module procTest_00_tb();

// geracao de clock e reset ---------------------------------------------------

reg clk, rst;

initial begin
    clk = 0;
    rst = 1;
    #1000.000000;
    rst = 0;
end

always #500.000000 clk = ~clk;

// instancia do processador ---------------------------------------------------

reg  signed [31:0] proc_io_in = 0;
wire signed [31:0] proc_io_out;
wire [0:0] proc_req_in;
wire [6:0] proc_out_en;

procTest_00 proc(clk,rst,proc_io_in,proc_io_out,proc_req_in,proc_out_en);

// portas de entrada ----------------------------------------------------------

// variaveis da porta 0
integer data_in_0;
reg signed [31:0] in_0 = 0;
reg req_in_0 = 0;

// abre um arquivo para leitura em cada porta
initial begin
    data_in_0 = $fopen("C:/Users/Ricardo/Documents/Dissertacao/banco_filtro/procTest_00/Simulation/input_0.txt", "r"); // coloque os seus dados de entrada neste arquivo
end

// decodifica portas de entrada
always @ (*) begin
    // decodificacao da porta 0
    if (proc_req_in == 1) proc_io_in = in_0;
    req_in_0 = proc_req_in == 1;
end

// implementa a leitura dos dados de entrada
integer scan_result;
always @ (negedge clk) begin  
    // lendo a porta 0
    if (data_in_0 != 0 && proc_req_in == 1) scan_result = $fscanf(data_in_0, "%d", in_0);
end

// portas de saida ------------------------------------------------------------

// variaveis da porta 1
integer data_out_1;
reg signed [31:0] out_sig_1 = 0;
reg out_en_1 = 0;

// variaveis da porta 2
integer data_out_2;
reg signed [31:0] out_sig_2 = 0;
reg out_en_2 = 0;

// variaveis da porta 3
integer data_out_3;
reg signed [31:0] out_sig_3 = 0;
reg out_en_3 = 0;

// variaveis da porta 4
integer data_out_4;
reg signed [31:0] out_sig_4 = 0;
reg out_en_4 = 0;

// variaveis da porta 5
integer data_out_5;
reg signed [31:0] out_sig_5 = 0;
reg out_en_5 = 0;

// variaveis da porta 6
integer data_out_6;
reg signed [31:0] out_sig_6 = 0;
reg out_en_6 = 0;

// abre um arquivo para escrita de cada porta
initial begin
    data_out_1 = $fopen("C:/Users/Ricardo/Documents/Dissertacao/banco_filtro/procTest_00/Simulation/output_1.txt", "w"); // veja os dados de saida neste arquivo
    data_out_2 = $fopen("C:/Users/Ricardo/Documents/Dissertacao/banco_filtro/procTest_00/Simulation/output_2.txt", "w"); // veja os dados de saida neste arquivo
    data_out_3 = $fopen("C:/Users/Ricardo/Documents/Dissertacao/banco_filtro/procTest_00/Simulation/output_3.txt", "w"); // veja os dados de saida neste arquivo
    data_out_4 = $fopen("C:/Users/Ricardo/Documents/Dissertacao/banco_filtro/procTest_00/Simulation/output_4.txt", "w"); // veja os dados de saida neste arquivo
    data_out_5 = $fopen("C:/Users/Ricardo/Documents/Dissertacao/banco_filtro/procTest_00/Simulation/output_5.txt", "w"); // veja os dados de saida neste arquivo
    data_out_6 = $fopen("C:/Users/Ricardo/Documents/Dissertacao/banco_filtro/procTest_00/Simulation/output_6.txt", "w"); // veja os dados de saida neste arquivo
end

// decodifica portas de saida
always @ (*) begin
    // decodificacao da porta 1
    if (proc_out_en == 2) out_sig_1 <= proc_io_out;
    out_en_1 = proc_out_en == 2;
    // decodificacao da porta 2
    if (proc_out_en == 4) out_sig_2 <= proc_io_out;
    out_en_2 = proc_out_en == 4;
    // decodificacao da porta 3
    if (proc_out_en == 8) out_sig_3 <= proc_io_out;
    out_en_3 = proc_out_en == 8;
    // decodificacao da porta 4
    if (proc_out_en == 16) out_sig_4 <= proc_io_out;
    out_en_4 = proc_out_en == 16;
    // decodificacao da porta 5
    if (proc_out_en == 32) out_sig_5 <= proc_io_out;
    out_en_5 = proc_out_en == 32;
    // decodificacao da porta 6
    if (proc_out_en == 64) out_sig_6 <= proc_io_out;
    out_en_6 = proc_out_en == 64;
end

// implementa escrita no arquivo
always @ (posedge clk) begin
    // escreve na porta 1
    if (out_en_1 == 1'b1) $fdisplay(data_out_1, "%0d", out_sig_1);
    // escreve na porta 2
    if (out_en_2 == 1'b1) $fdisplay(data_out_2, "%0d", out_sig_2);
    // escreve na porta 3
    if (out_en_3 == 1'b1) $fdisplay(data_out_3, "%0d", out_sig_3);
    // escreve na porta 4
    if (out_en_4 == 1'b1) $fdisplay(data_out_4, "%0d", out_sig_4);
    // escreve na porta 5
    if (out_en_5 == 1'b1) $fdisplay(data_out_5, "%0d", out_sig_5);
    // escreve na porta 6
    if (out_en_6 == 1'b1) $fdisplay(data_out_6, "%0d", out_sig_6);
end

// cadastro de sinais, barra de progresso e finish ----------------------------

integer progress, chrys;
initial begin

    $dumpfile("procTest_00_tb.vcd");

    $dumpvars(0,procTest_00_tb.clk);
    $dumpvars(0,procTest_00_tb.rst);
    $dumpvars(0,procTest_00_tb.proc.req_in_sim_0);
    $dumpvars(0,procTest_00_tb.proc.in_sim_0);
    $dumpvars(0,procTest_00_tb.proc.out_en_sim_1);
    $dumpvars(0,procTest_00_tb.proc.out_sig_1);
    $dumpvars(0,procTest_00_tb.proc.out_en_sim_2);
    $dumpvars(0,procTest_00_tb.proc.out_sig_2);
    $dumpvars(0,procTest_00_tb.proc.out_en_sim_3);
    $dumpvars(0,procTest_00_tb.proc.out_sig_3);
    $dumpvars(0,procTest_00_tb.proc.out_en_sim_4);
    $dumpvars(0,procTest_00_tb.proc.out_sig_4);
    $dumpvars(0,procTest_00_tb.proc.out_en_sim_5);
    $dumpvars(0,procTest_00_tb.proc.out_sig_5);
    $dumpvars(0,procTest_00_tb.proc.out_en_sim_6);
    $dumpvars(0,procTest_00_tb.proc.out_sig_6);
    $dumpvars(0,procTest_00_tb.proc.valr2);
    $dumpvars(0,procTest_00_tb.proc.linetabs);
    $dumpvars(0,procTest_00_tb.proc.me1_f_ifft_v_N_e_);
    $dumpvars(0,procTest_00_tb.proc.me1_f_ifft_v_mmax_e_);
    $dumpvars(0,procTest_00_tb.proc.me1_f_ifft_v_istep_e_);
    $dumpvars(0,procTest_00_tb.proc.me1_f_ifft_v_m_e_);
    $dumpvars(0,procTest_00_tb.proc.me1_f_ifft_v_ind_e_);
    $dumpvars(0,procTest_00_tb.proc.me1_f_ifft_v_sind_e_);
    $dumpvars(0,procTest_00_tb.proc.me1_f_ifft_v_k_e_);
    $dumpvars(0,procTest_00_tb.proc.me1_f_ifft_v_j_e_);
    $dumpvars(0,procTest_00_tb.proc.comp_me3_f_ifft_v_temp_e_);
    $dumpvars(0,procTest_00_tb.proc.me1_f_main_v_sample_count_e_);
    $dumpvars(0,procTest_00_tb.proc.me1_f_main_v_output_count_e_);
    $dumpvars(0,procTest_00_tb.proc.me1_f_main_v_M_e_);
    $dumpvars(0,procTest_00_tb.proc.me1_f_main_v_fft_limit_e_);
    $dumpvars(0,procTest_00_tb.proc.me1_f_main_v_k_e_);
    $dumpvars(0,procTest_00_tb.proc.me1_f_main_v_mm_e_);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0000);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0001);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0002);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0003);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0004);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0005);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0006);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0007);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0008);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0009);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0010);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0011);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0012);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0013);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0014);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0015);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0016);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0017);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0018);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0019);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0020);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0021);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0022);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0023);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0024);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0025);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0026);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0027);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0028);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0029);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0030);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0031);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0032);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0033);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0034);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0035);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0036);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0037);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0038);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0039);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0040);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0041);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0042);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0043);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0044);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0045);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0046);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0047);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0048);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0049);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0050);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0051);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0052);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0053);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0054);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0055);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0056);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0057);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0058);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0059);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0060);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0061);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0062);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0063);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0064);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0065);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0066);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0067);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0068);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0069);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0070);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0071);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0072);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0073);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0074);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0075);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0076);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0077);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0078);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0079);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0080);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0081);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0082);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0083);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0084);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0085);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0086);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0087);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0088);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0089);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0090);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0091);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0092);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0093);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0094);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0095);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0096);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0097);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0098);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0099);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0100);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0101);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0102);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0103);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0104);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0105);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0106);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0107);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0108);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0109);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0110);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0111);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0112);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0113);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0114);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0115);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0116);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0117);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0118);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0119);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0120);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0121);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0122);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0123);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0124);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0125);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0126);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0127);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0128);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0129);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0130);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0131);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0132);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0133);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0134);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0135);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0136);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0137);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0138);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0139);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0140);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0141);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0142);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0143);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0144);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0145);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0146);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0147);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0148);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0149);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0150);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0151);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0152);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0153);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0154);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0155);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0156);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0157);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0158);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0159);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0160);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0161);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0162);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0163);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0164);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0165);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0166);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0167);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0168);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0169);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0170);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0171);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0172);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0173);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0174);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0175);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0176);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0177);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0178);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0179);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0180);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0181);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0182);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0183);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0184);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0185);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0186);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0187);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0188);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0189);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0190);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0191);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0192);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0193);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0194);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0195);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0196);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0197);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0198);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0199);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0200);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0201);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0202);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0203);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0204);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0205);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0206);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0207);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0208);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0209);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0210);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0211);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0212);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0213);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0214);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0215);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0216);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0217);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0218);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0219);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0220);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0221);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0222);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0223);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0224);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0225);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0226);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0227);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0228);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0229);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0230);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0231);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0232);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0233);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0234);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0235);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0236);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0237);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0238);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0239);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0240);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0241);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0242);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0243);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0244);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0245);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0246);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0247);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0248);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0249);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0250);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0251);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0252);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0253);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0254);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_E0_e_0255);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0000);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0001);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0002);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0003);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0004);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0005);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0006);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0007);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0008);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0009);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0010);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0011);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0012);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0013);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0014);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0015);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0016);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0017);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0018);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0019);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0020);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0021);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0022);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0023);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0024);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0025);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0026);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0027);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0028);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0029);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0030);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0031);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0032);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0033);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0034);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0035);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0036);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0037);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0038);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0039);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0040);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0041);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0042);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0043);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0044);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0045);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0046);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0047);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0048);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0049);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0050);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0051);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0052);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0053);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0054);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0055);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0056);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0057);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0058);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0059);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0060);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0061);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0062);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0063);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0064);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0065);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0066);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0067);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0068);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0069);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0070);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0071);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0072);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0073);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0074);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0075);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0076);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0077);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0078);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0079);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0080);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0081);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0082);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0083);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0084);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0085);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0086);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0087);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0088);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0089);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0090);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0091);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0092);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0093);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0094);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0095);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0096);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0097);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0098);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0099);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0100);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0101);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0102);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0103);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0104);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0105);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0106);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0107);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0108);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0109);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0110);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0111);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0112);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0113);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0114);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0115);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0116);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0117);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0118);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0119);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0120);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0121);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0122);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0123);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0124);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0125);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0126);
    $dumpvars(0,procTest_00_tb.proc.comp_arr_me3_f_global_v_wpv_e_0127);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0000);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0001);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0002);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0003);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0004);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0005);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0006);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0007);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0008);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0009);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0010);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0011);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0012);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0013);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0014);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0015);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0016);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0017);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0018);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0019);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0020);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0021);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0022);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0023);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0024);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0025);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0026);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0027);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0028);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0029);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0030);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0031);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0032);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0033);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0034);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0035);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0036);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0037);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0038);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0039);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0040);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0041);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0042);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0043);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0044);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0045);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0046);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0047);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0048);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0049);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0050);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0051);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0052);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0053);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0054);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0055);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0056);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0057);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0058);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0059);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0060);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0061);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0062);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0063);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0064);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0065);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0066);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0067);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0068);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0069);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0070);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0071);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0072);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0073);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0074);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0075);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0076);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0077);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0078);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0079);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0080);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0081);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0082);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0083);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0084);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0085);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0086);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0087);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0088);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0089);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0090);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0091);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0092);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0093);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0094);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0095);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0096);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0097);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0098);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0099);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0100);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0101);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0102);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0103);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0104);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0105);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0106);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0107);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0108);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0109);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0110);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0111);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0112);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0113);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0114);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0115);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0116);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0117);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0118);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0119);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0120);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0121);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0122);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0123);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0124);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0125);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0126);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0127);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0128);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0129);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0130);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0131);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0132);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0133);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0134);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0135);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0136);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0137);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0138);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0139);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0140);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0141);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0142);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0143);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0144);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0145);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0146);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0147);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0148);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0149);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0150);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0151);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0152);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0153);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0154);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0155);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0156);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0157);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0158);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0159);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0160);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0161);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0162);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0163);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0164);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0165);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0166);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0167);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0168);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0169);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0170);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0171);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0172);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0173);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0174);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0175);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0176);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0177);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0178);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0179);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0180);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0181);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0182);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0183);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0184);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0185);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0186);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0187);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0188);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0189);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0190);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0191);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0192);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0193);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0194);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0195);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0196);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0197);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0198);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0199);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0200);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0201);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0202);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0203);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0204);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0205);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0206);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0207);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0208);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0209);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0210);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0211);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0212);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0213);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0214);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0215);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0216);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0217);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0218);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0219);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0220);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0221);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0222);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0223);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0224);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0225);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0226);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0227);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0228);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0229);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0230);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0231);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0232);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0233);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0234);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0235);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0236);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0237);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0238);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0239);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0240);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0241);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0242);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0243);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0244);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0245);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0246);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0247);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0248);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0249);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0250);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0251);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0252);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0253);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0254);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_real_e_0255);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0000);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0001);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0002);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0003);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0004);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0005);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0006);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0007);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0008);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0009);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0010);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0011);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0012);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0013);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0014);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0015);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0016);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0017);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0018);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0019);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0020);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0021);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0022);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0023);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0024);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0025);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0026);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0027);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0028);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0029);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0030);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0031);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0032);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0033);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0034);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0035);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0036);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0037);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0038);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0039);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0040);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0041);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0042);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0043);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0044);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0045);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0046);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0047);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0048);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0049);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0050);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0051);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0052);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0053);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0054);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0055);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0056);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0057);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0058);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0059);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0060);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0061);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0062);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0063);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0064);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0065);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0066);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0067);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0068);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0069);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0070);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0071);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0072);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0073);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0074);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0075);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0076);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0077);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0078);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0079);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0080);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0081);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0082);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0083);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0084);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0085);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0086);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0087);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0088);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0089);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0090);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0091);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0092);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0093);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0094);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0095);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0096);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0097);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0098);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0099);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0100);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0101);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0102);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0103);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0104);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0105);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0106);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0107);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0108);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0109);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0110);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0111);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0112);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0113);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0114);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0115);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0116);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0117);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0118);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0119);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0120);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0121);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0122);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0123);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0124);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0125);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0126);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0127);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0128);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0129);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0130);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0131);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0132);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0133);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0134);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0135);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0136);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0137);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0138);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0139);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0140);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0141);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0142);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0143);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0144);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0145);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0146);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0147);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0148);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0149);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0150);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0151);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0152);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0153);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0154);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0155);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0156);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0157);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0158);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0159);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0160);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0161);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0162);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0163);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0164);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0165);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0166);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0167);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0168);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0169);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0170);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0171);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0172);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0173);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0174);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0175);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0176);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0177);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0178);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0179);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0180);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0181);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0182);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0183);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0184);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0185);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0186);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0187);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0188);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0189);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0190);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0191);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0192);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0193);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0194);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0195);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0196);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0197);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0198);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0199);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0200);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0201);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0202);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0203);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0204);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0205);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0206);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0207);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0208);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0209);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0210);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0211);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0212);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0213);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0214);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0215);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0216);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0217);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0218);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0219);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0220);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0221);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0222);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0223);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0224);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0225);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0226);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0227);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0228);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0229);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0230);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0231);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0232);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0233);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0234);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0235);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0236);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0237);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0238);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0239);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0240);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0241);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0242);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0243);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0244);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0245);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0246);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0247);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0248);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0249);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0250);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0251);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0252);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0253);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0254);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_output_buffer_imag_e_0255);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0000);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0001);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0002);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0003);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0004);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0005);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0006);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0007);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0008);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0009);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0010);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0011);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0012);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0013);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0014);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0015);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0016);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0017);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0018);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0019);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0020);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0021);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0022);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0023);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0024);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0025);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0026);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0027);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0028);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0029);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0030);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0031);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0032);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0033);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0034);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0035);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0036);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0037);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0038);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0039);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0040);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0041);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0042);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0043);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0044);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0045);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0046);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0047);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0048);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0049);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0050);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0051);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0052);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0053);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0054);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0055);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0056);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0057);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0058);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0059);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0060);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0061);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0062);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0063);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0064);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0065);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0066);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0067);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0068);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0069);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0070);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0071);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0072);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0073);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0074);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0075);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0076);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0077);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0078);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0079);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0080);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0081);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0082);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0083);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0084);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0085);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0086);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0087);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0088);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0089);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0090);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0091);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0092);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0093);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0094);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0095);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0096);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0097);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0098);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0099);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0100);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0101);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0102);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0103);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0104);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0105);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0106);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0107);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0108);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0109);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0110);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0111);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0112);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0113);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0114);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0115);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0116);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0117);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0118);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0119);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0120);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0121);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0122);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0123);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0124);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0125);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0126);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0127);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0128);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0129);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0130);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0131);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0132);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0133);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0134);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0135);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0136);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0137);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0138);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0139);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0140);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0141);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0142);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0143);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0144);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0145);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0146);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0147);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0148);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0149);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0150);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0151);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0152);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0153);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0154);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0155);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0156);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0157);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0158);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0159);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0160);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0161);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0162);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0163);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0164);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0165);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0166);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0167);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0168);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0169);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0170);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0171);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0172);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0173);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0174);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0175);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0176);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0177);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0178);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0179);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0180);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0181);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0182);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0183);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0184);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0185);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0186);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0187);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0188);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0189);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0190);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0191);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0192);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0193);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0194);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0195);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0196);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0197);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0198);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0199);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0200);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0201);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0202);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0203);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0204);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0205);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0206);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0207);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0208);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0209);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0210);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0211);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0212);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0213);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0214);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0215);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0216);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0217);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0218);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0219);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0220);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0221);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0222);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0223);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0224);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0225);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0226);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0227);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0228);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0229);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0230);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0231);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0232);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0233);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0234);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0235);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0236);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0237);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0238);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0239);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0240);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0241);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0242);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0243);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0244);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0245);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0246);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0247);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0248);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0249);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0250);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0251);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0252);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0253);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0254);
    $dumpvars(0,procTest_00_tb.proc.arr_me2_f_main_v_buffer_e_0255);
    $dumpvars(0,procTest_00_tb.proc.p_procTest_00.core.instr_fetch.genblk2.isp.pointeri);
    $dumpvars(0,procTest_00_tb.proc.p_procTest_00.core.instr_fetch.genblk2.isp.fl_max);
    $dumpvars(0,procTest_00_tb.proc.p_procTest_00.core.instr_fetch.genblk2.isp.fl_full);
    $dumpvars(0,procTest_00_tb.proc.p_procTest_00.core.sp.pointeri);
    $dumpvars(0,procTest_00_tb.proc.p_procTest_00.core.sp.fl_max);
    $dumpvars(0,procTest_00_tb.proc.p_procTest_00.core.sp.fl_full);
    $dumpvars(0,procTest_00_tb.proc.p_procTest_00.core.ula.delta_float);
    $dumpvars(0,procTest_00_tb.proc.p_procTest_00.core.ula.delta_int);

    progress = $fopen("progress.txt", "w");
    for (chrys = 10; chrys <= 100; chrys = chrys + 10) begin
        #800000000.000000;
        $fdisplay(progress,"%0d",chrys);
        $fflush(progress);
    end

    $fclose(progress);
    $finish;

end

endmodule
